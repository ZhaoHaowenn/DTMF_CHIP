// Created on Wed Mar 15 17:09:43 2006
module accum_stat (
	accum,
	ar,
	bio,
	gez,
	gz,
	nz,
	z,
	lz,
	lez,
	ov,
	arnz,
	bioz );
   input [32:0] accum;
   input [15:0] ar;
   input bio;
   output gez;
   output gz;
   output nz;
   output z;
   output lz;
   output lez;
   input ov;
   output arnz;
   output bioz;

   // Internal wires
   wire n_6309;
   wire n_73;
   wire n_46;
   wire n_49;
   wire n_53;
   wire n_56;
   wire n_58;
   wire n_61;
   wire n_64;
   wire n_68;
   wire n_71;
   wire n_76;
   wire n_79;
   wire n_83;
   wire n_87;

   INVXL i_9530 ( .Y (lz),
	.A (n_6309) );
   INVXL i_9529 ( .Y (n_6309),
	.A (accum[31]) );
   NOR2X1 i_4403 ( .Y (gz),
	.B (n_73),
	.A (lz) );
   NOR4X1 i_43 ( .Y (n_46),
	.D (accum[1]),
	.C (accum[0]),
	.B (accum[3]),
	.A (accum[2]) );
   NOR4X1 i_40 ( .Y (n_49),
	.D (accum[5]),
	.C (accum[4]),
	.B (accum[7]),
	.A (accum[6]) );
   NOR4X1 i_36 ( .Y (n_53),
	.D (accum[9]),
	.C (accum[8]),
	.B (accum[11]),
	.A (accum[10]) );
   NOR4X1 i_33 ( .Y (n_56),
	.D (accum[13]),
	.C (accum[12]),
	.B (accum[15]),
	.A (accum[14]) );
   NAND4X1 i_45 ( .Y (n_58),
	.D (n_46),
	.C (n_49),
	.B (n_53),
	.A (n_56) );
   OR4X1 i_28 ( .Y (n_61),
	.D (accum[17]),
	.C (accum[16]),
	.B (accum[19]),
	.A (accum[18]) );
   NOR4X1 i_25 ( .Y (n_64),
	.D (accum[21]),
	.C (accum[20]),
	.B (accum[23]),
	.A (accum[22]) );
   OR4X1 i_21 ( .Y (n_68),
	.D (accum[25]),
	.C (accum[24]),
	.B (accum[27]),
	.A (accum[26]) );
   OR4X1 i_22 ( .Y (n_71),
	.D (n_68),
	.C (accum[30]),
	.B (accum[29]),
	.A (accum[28]) );
   NOR4BX1 i_09004 ( .Y (n_73),
	.D (n_71),
	.C (n_61),
	.B (n_58),
	.AN (n_64) );
   NOR4X1 i_13 ( .Y (n_76),
	.D (ar[1]),
	.C (ar[0]),
	.B (ar[3]),
	.A (ar[2]) );
   NOR4X1 i_10 ( .Y (n_79),
	.D (ar[5]),
	.C (ar[4]),
	.B (ar[7]),
	.A (ar[6]) );
   NOR4X1 i_6 ( .Y (n_83),
	.D (ar[9]),
	.C (ar[8]),
	.B (ar[11]),
	.A (ar[10]) );
   NOR4X1 i_3 ( .Y (n_87),
	.D (ar[13]),
	.C (ar[12]),
	.B (ar[15]),
	.A (ar[14]) );
   OAI21XL i_4401 ( .Y (gez),
	.B0 (nz),
	.A1 (n_73),
	.A0 (lz) );
   NAND2BX1 i_4406 ( .Y (nz),
	.B (n_73),
	.AN (lz) );
   OR2X1 i_4405 ( .Y (lez),
	.B (n_73),
	.A (lz) );
   NAND4X1 i_342308 ( .Y (arnz),
	.D (n_76),
	.C (n_79),
	.B (n_83),
	.A (n_87) );
   INVX1 i_3339 ( .Y (bioz),
	.A (bio) );
endmodule

module alu_32 (
	ovm,
	op_a,
	op_b,
	result,
	cmd );
   input ovm;
   input [31:0] op_a;
   input [31:0] op_b;
   output [32:0] result;
   input [3:0] cmd;

   // Internal wires
   wire n_2382;
   wire n_911;
   wire n_1618;
   wire n_1830;
   wire n_1831;
   wire n_1827;
   wire n_1616;
   wire n_1617;
   wire n_906;
   wire n_1880;
   wire n_1936;
   wire n_1614;
   wire n_949;
   wire n_3062;
   wire n_1613;
   wire n_879;
   wire n_1611;
   wire n_1754;
   wire n_1612;
   wire n_1806;
   wire n_1758;
   wire n_946;
   wire n_1609;
   wire n_907;
   wire n_3060;
   wire n_1598;
   wire n_2360;
   wire n_1727;
   wire n_2378;
   wire n_2370;
   wire n_1699;
   wire n_1596;
   wire n_1600;
   wire n_2372;
   wire n_1589;
   wire n_1599;
   wire n_1708;
   wire n_1716;
   wire n_2264;
   wire n_2300;
   wire n_2299;
   wire n_1593;
   wire n_1594;
   wire n_1441;
   wire n_1395;
   wire n_1494;
   wire n_1592;
   wire n_2295;
   wire n_2259;
   wire n_2294;
   wire n_1586;
   wire n_1587;
   wire n_2260;
   wire n_1485;
   wire n_925;
   wire n_1487;
   wire n_1585;
   wire n_1582;
   wire n_1571;
   wire n_2341;
   wire n_2358;
   wire n_1573;
   wire n_3095;
   wire n_1579;
   wire n_1566;
   wire n_2346;
   wire n_2349;
   wire n_1568;
   wire n_2285;
   wire n_2351;
   wire n_1563;
   wire n_1572;
   wire n_2344;
   wire n_1738;
   wire n_1835;
   wire n_1879;
   wire n_1565;
   wire n_1567;
   wire n_1881;
   wire n_1390;
   wire n_1467;
   wire n_1762;
   wire n_1757;
   wire n_1559;
   wire n_1561;
   wire n_1462;
   wire n_927;
   wire n_1383;
   wire n_1557;
   wire n_1546;
   wire n_2323;
   wire n_2339;
   wire n_2333;
   wire n_1647;
   wire n_1543;
   wire n_1548;
   wire n_1907;
   wire n_1536;
   wire n_1547;
   wire n_1637;
   wire n_1544;
   wire n_2233;
   wire n_2265;
   wire n_1540;
   wire n_1541;
   wire n_2234;
   wire n_1443;
   wire n_1539;
   wire n_2228;
   wire n_1533;
   wire n_1534;
   wire n_1436;
   wire n_929;
   wire n_1532;
   wire n_1529;
   wire n_1518;
   wire n_2313;
   wire n_2321;
   wire n_2315;
   wire n_1516;
   wire n_1520;
   wire n_1930;
   wire n_1932;
   wire n_1513;
   wire n_1519;
   wire n_1510;
   wire n_1499;
   wire n_2293;
   wire n_2311;
   wire n_2303;
   wire n_1496;
   wire n_1501;
   wire n_2305;
   wire n_1500;
   wire n_1497;
   wire n_2198;
   wire n_1493;
   wire n_1339;
   wire n_1297;
   wire n_1392;
   wire n_1492;
   wire n_2229;
   wire n_2193;
   wire n_1486;
   wire n_2194;
   wire n_1385;
   wire n_1482;
   wire n_1471;
   wire n_2276;
   wire n_2291;
   wire n_2282;
   wire n_1469;
   wire n_1473;
   wire n_1464;
   wire n_1472;
   wire n_1843;
   wire n_1877;
   wire n_1838;
   wire n_1466;
   wire n_1293;
   wire n_1365;
   wire n_1804;
   wire n_1770;
   wire n_1765;
   wire n_1461;
   wire n_1360;
   wire n_931;
   wire n_1286;
   wire n_1459;
   wire n_1448;
   wire n_2258;
   wire n_2274;
   wire n_2268;
   wire n_1445;
   wire n_1450;
   wire n_1903;
   wire n_1449;
   wire n_1446;
   wire n_2167;
   wire n_2199;
   wire n_1442;
   wire n_2168;
   wire n_1340;
   wire n_2162;
   wire n_1435;
   wire n_1334;
   wire n_933;
   wire n_1434;
   wire n_1431;
   wire n_1420;
   wire n_2248;
   wire n_2256;
   wire n_2250;
   wire n_1418;
   wire n_1422;
   wire n_1413;
   wire n_1421;
   wire n_1846;
   wire n_1847;
   wire n_1415;
   wire n_1416;
   wire n_1875;
   wire n_903;
   wire n_1773;
   wire n_1774;
   wire n_1410;
   wire n_1411;
   wire n_1802;
   wire n_943;
   wire n_1408;
   wire n_1397;
   wire n_2227;
   wire n_2246;
   wire n_2237;
   wire n_1394;
   wire n_1399;
   wire n_2174;
   wire n_2239;
   wire n_1387;
   wire n_1398;
   wire n_2132;
   wire n_1391;
   wire n_1244;
   wire n_1198;
   wire n_1294;
   wire n_2163;
   wire n_2127;
   wire n_1384;
   wire n_2128;
   wire n_1287;
   wire n_1380;
   wire n_1369;
   wire n_2210;
   wire n_2225;
   wire n_2216;
   wire n_1367;
   wire n_1371;
   wire n_2153;
   wire n_2218;
   wire n_1362;
   wire n_1370;
   wire n_1851;
   wire n_1364;
   wire n_1193;
   wire n_1268;
   wire n_1778;
   wire n_1359;
   wire n_1264;
   wire n_935;
   wire n_1186;
   wire n_1357;
   wire n_1346;
   wire n_2192;
   wire n_2208;
   wire n_2202;
   wire n_1343;
   wire n_1348;
   wire n_1899;
   wire n_1337;
   wire n_1347;
   wire n_1344;
   wire n_2103;
   wire n_1245;
   wire n_1341;
   wire n_2102;
   wire n_2133;
   wire n_2097;
   wire n_1333;
   wire n_1238;
   wire n_937;
   wire n_1332;
   wire n_1329;
   wire n_1318;
   wire n_2182;
   wire n_2190;
   wire n_2184;
   wire n_1316;
   wire n_1320;
   wire n_1924;
   wire n_1926;
   wire n_1314;
   wire n_1319;
   wire n_1310;
   wire n_1299;
   wire n_2161;
   wire n_2180;
   wire n_2171;
   wire n_1296;
   wire n_1301;
   wire n_1291;
   wire n_1300;
   wire n_2066;
   wire n_855;
   wire n_1187;
   wire n_2062;
   wire n_1288;
   wire n_2098;
   wire n_2061;
   wire n_1283;
   wire n_1272;
   wire n_2144;
   wire n_2159;
   wire n_2150;
   wire n_1270;
   wire n_1274;
   wire n_1267;
   wire n_1273;
   wire n_1873;
   wire n_1863;
   wire n_1167;
   wire n_3092;
   wire n_1800;
   wire n_1790;
   wire n_1162;
   wire n_2080;
   wire n_1262;
   wire n_1251;
   wire n_2126;
   wire n_2142;
   wire n_2136;
   wire n_1248;
   wire n_1253;
   wire n_1895;
   wire n_1252;
   wire n_1249;
   wire n_2039;
   wire n_1144;
   wire n_1100;
   wire n_2004;
   wire n_1246;
   wire n_2038;
   wire n_2067;
   wire n_1090;
   wire n_1137;
   wire n_942;
   wire n_1239;
   wire n_862;
   wire n_1237;
   wire n_1234;
   wire n_1223;
   wire n_2116;
   wire n_2124;
   wire n_2118;
   wire n_1221;
   wire n_1225;
   wire n_1217;
   wire n_1224;
   wire n_1053;
   wire n_1097;
   wire n_1870;
   wire n_1219;
   wire n_1862;
   wire n_1859;
   wire n_1218;
   wire n_1797;
   wire n_1799;
   wire n_861;
   wire n_1786;
   wire n_1213;
   wire n_1211;
   wire n_1200;
   wire n_2096;
   wire n_2114;
   wire n_2106;
   wire n_1197;
   wire n_1202;
   wire n_2108;
   wire n_1191;
   wire n_1201;
   wire n_2003;
   wire n_1976;
   wire n_3089;
   wire n_1194;
   wire n_1997;
   wire n_1972;
   wire n_1188;
   wire n_1089;
   wire n_1785;
   wire n_860;
   wire n_1183;
   wire n_1172;
   wire n_2079;
   wire n_2094;
   wire n_2085;
   wire n_1170;
   wire n_1174;
   wire n_2017;
   wire n_2087;
   wire n_1166;
   wire n_1173;
   wire n_1869;
   wire n_3085;
   wire n_1871;
   wire n_1168;
   wire n_2020;
   wire n_1798;
   wire n_857;
   wire n_2013;
   wire n_1160;
   wire n_1149;
   wire n_2060;
   wire n_2077;
   wire n_2070;
   wire n_1146;
   wire n_1151;
   wire n_1891;
   wire n_1150;
   wire n_1147;
   wire n_856;
   wire n_1998;
   wire n_1136;
   wire n_1135;
   wire n_1132;
   wire n_1122;
   wire n_2049;
   wire n_2059;
   wire n_1915;
   wire n_2052;
   wire n_1917;
   wire n_1129;
   wire n_2053;
   wire n_1119;
   wire n_1123;
   wire n_3076;
   wire n_2051;
   wire n_1116;
   wire n_1113;
   wire n_1103;
   wire n_2028;
   wire n_2048;
   wire n_2037;
   wire n_1110;
   wire n_2042;
   wire n_1099;
   wire n_1104;
   wire n_1096;
   wire n_1095;
   wire n_2036;
   wire n_1092;
   wire n_1787;
   wire n_1087;
   wire n_1085;
   wire n_1084;
   wire n_2025;
   wire n_1076;
   wire n_2019;
   wire n_2021;
   wire n_1073;
   wire n_1078;
   wire n_1071;
   wire n_1072;
   wire n_2018;
   wire n_1070;
   wire n_1068;
   wire n_1066;
   wire n_1056;
   wire n_1995;
   wire n_2011;
   wire n_2001;
   wire n_1063;
   wire n_2005;
   wire n_1052;
   wire n_1057;
   wire n_2000;
   wire n_1048;
   wire n_1045;
   wire n_1042;
   wire n_1032;
   wire n_1984;
   wire n_1994;
   wire n_1987;
   wire n_1039;
   wire n_1988;
   wire n_1029;
   wire n_1033;
   wire n_1986;
   wire n_1026;
   wire n_1023;
   wire n_1013;
   wire n_1970;
   wire n_1983;
   wire n_1975;
   wire n_1020;
   wire n_1977;
   wire n_1014;
   wire n_1974;
   wire n_1006;
   wire n_1002;
   wire n_992;
   wire n_1959;
   wire n_1969;
   wire n_1962;
   wire n_999;
   wire n_3083;
   wire n_988;
   wire n_993;
   wire n_1795;
   wire n_1961;
   wire n_986;
   wire n_983;
   wire n_9076575;
   wire n_827;
   wire n_984;
   wire n_981;
   wire n_1957;
   wire n_976;
   wire n_1946;
   wire n_974;
   wire n_978;
   wire n_973;
   wire n_1955;
   wire n_1950;
   wire n_1733;
   wire n_971;
   wire n_970;
   wire n_1938;
   wire n_1918;
   wire n_967;
   wire n_1810;
   wire n_1883;
   wire n_868;
   wire n_964;
   wire n_958;
   wire n_1944;
   wire n_1942;
   wire n_963;
   wire n_962;
   wire n_951;
   wire n_1713;
   wire n_885;
   wire n_955;
   wire n_954;
   wire n_952;
   wire n_1743;
   wire n_3070;
   wire n_1809;
   wire n_1751;
   wire n_1766;
   wire n_945;
   wire n_1782;
   wire n_944;
   wire n_1781;
   wire n_940;
   wire n_923;
   wire n_921;
   wire n_913;
   wire n_1703;
   wire n_1812;
   wire n_917;
   wire n_915;
   wire n_1816;
   wire n_3086;
   wire n_1815;
   wire n_1822;
   wire n_1823;
   wire n_1819;
   wire n_909;
   wire n_1882;
   wire n_1839;
   wire n_905;
   wire n_904;
   wire n_1854;
   wire n_1855;
   wire n_2324;
   wire n_2362;
   wire n_882;
   wire n_2029;
   wire n_1789;
   wire n_3087;
   wire n_3065;
   wire n_828;
   wire n_1640;
   wire n_3069;
   wire n_1620;
   wire n_1622;
   wire n_1623;
   wire n_1630;
   wire n_2387;
   wire n_1632;
   wire n_2325;
   wire n_1635;
   wire n_2361;
   wire n_1639;
   wire n_1645;
   wire n_2367;
   wire n_1646;
   wire n_2330;
   wire n_2329;
   wire n_2366;
   wire n_1648;
   wire n_1650;
   wire n_2402;
   wire n_2401;
   wire n_1652;
   wire n_2390;
   wire n_1654;
   wire n_1653;
   wire n_2393;
   wire n_1911;
   wire n_1655;
   wire n_1656;
   wire n_3068;
   wire n_1661;
   wire n_2397;
   wire n_2404;
   wire n_1665;
   wire n_2408;
   wire n_1670;
   wire n_2417;
   wire n_1672;
   wire n_1674;
   wire n_2411;
   wire n_3077;
   wire n_1676;
   wire n_2413;
   wire n_1678;
   wire n_2409;
   wire n_1681;
   wire n_1682;
   wire n_1683;
   wire n_2406;
   wire n_1689;
   wire n_2423;
   wire n_1692;
   wire n_1696;
   wire n_1697;
   wire n_1700;
   wire n_1698;
   wire n_2399;
   wire n_3066;
   wire n_1704;
   wire n_1705;
   wire n_1706;
   wire n_1709;
   wire n_1710;
   wire n_2391;
   wire n_2426;
   wire n_1714;
   wire n_1736;
   wire n_2434;
   wire n_2436;
   wire n_1720;
   wire n_2431;
   wire n_3088;
   wire n_1722;
   wire n_1723;
   wire n_2425;
   wire n_2441;
   wire n_1730;
   wire n_1740;
   wire n_1949;
   wire n_1734;
   wire n_1741;
   wire n_1742;
   wire n_1744;
   wire n_1745;
   wire n_1746;
   wire n_1747;
   wire n_1748;
   wire n_1749;
   wire n_1750;
   wire n_1752;
   wire n_1753;
   wire n_1755;
   wire n_1756;
   wire n_1760;
   wire n_1761;
   wire n_1763;
   wire n_1764;
   wire n_1768;
   wire n_1769;
   wire n_1771;
   wire n_1772;
   wire n_1776;
   wire n_1777;
   wire n_1779;
   wire n_1780;
   wire n_1784;
   wire n_3074;
   wire n_1788;
   wire n_1792;
   wire n_1793;
   wire n_1794;
   wire n_1808;
   wire n_1813;
   wire n_1814;
   wire n_1817;
   wire n_1818;
   wire n_1820;
   wire n_1821;
   wire n_1825;
   wire n_1826;
   wire n_1828;
   wire n_1829;
   wire n_1833;
   wire n_1834;
   wire n_1836;
   wire n_1837;
   wire n_1841;
   wire n_1842;
   wire n_1844;
   wire n_1845;
   wire n_1849;
   wire n_1850;
   wire n_1852;
   wire n_1853;
   wire n_1857;
   wire n_1858;
   wire n_1860;
   wire n_1861;
   wire n_1865;
   wire n_1866;
   wire n_1867;
   wire n_1868;
   wire n_1885;
   wire n_1886;
   wire n_1887;
   wire n_1888;
   wire n_1892;
   wire n_1893;
   wire n_1896;
   wire n_1900;
   wire n_1901;
   wire n_1904;
   wire n_1905;
   wire n_1908;
   wire n_1909;
   wire n_1912;
   wire n_166;
   wire n_1919;
   wire n_1921;
   wire n_1927;
   wire n_1933;
   wire n_1947;
   wire n_3075;
   wire n_3063;
   wire n_1965;
   wire n_1966;
   wire n_1968;
   wire n_1971;
   wire n_3084;
   wire n_1979;
   wire n_1980;
   wire n_1982;
   wire n_3067;
   wire n_3081;
   wire n_1990;
   wire n_1991;
   wire n_1993;
   wire n_1996;
   wire n_2002;
   wire n_3082;
   wire n_2007;
   wire n_2008;
   wire n_2010;
   wire n_2016;
   wire n_3079;
   wire n_2023;
   wire n_2035;
   wire n_2040;
   wire n_3080;
   wire n_2044;
   wire n_2045;
   wire n_2047;
   wire n_3078;
   wire n_2055;
   wire n_2056;
   wire n_2058;
   wire n_2071;
   wire n_2072;
   wire n_2074;
   wire n_2076;
   wire n_3073;
   wire n_2083;
   wire n_2088;
   wire n_2089;
   wire n_2091;
   wire n_2093;
   wire n_2109;
   wire n_2111;
   wire n_2113;
   wire n_2119;
   wire n_2121;
   wire n_2123;
   wire n_2137;
   wire n_2139;
   wire n_2141;
   wire n_2154;
   wire n_2156;
   wire n_2158;
   wire n_2175;
   wire n_2177;
   wire n_2179;
   wire n_2185;
   wire n_2187;
   wire n_2189;
   wire n_2203;
   wire n_2205;
   wire n_2207;
   wire n_2219;
   wire n_2220;
   wire n_2222;
   wire n_2224;
   wire n_2241;
   wire n_2243;
   wire n_2245;
   wire n_2251;
   wire n_2253;
   wire n_2255;
   wire n_2269;
   wire n_2271;
   wire n_2273;
   wire n_2286;
   wire n_2288;
   wire n_2290;
   wire n_2306;
   wire n_2308;
   wire n_2310;
   wire n_2316;
   wire n_2318;
   wire n_2320;
   wire n_2334;
   wire n_2336;
   wire n_2338;
   wire n_2342;
   wire n_3071;
   wire n_2352;
   wire n_2353;
   wire n_2355;
   wire n_2357;
   wire n_3093;
   wire n_2373;
   wire n_2375;
   wire n_2377;
   wire n_2383;
   wire n_2384;
   wire n_2385;
   wire n_2394;
   wire n_3064;
   wire n_2395;
   wire n_3090;
   wire n_3091;
   wire n_2418;
   wire n_2420;
   wire n_2422;
   wire n_2428;
   wire n_2437;
   wire n_2439;

   NOR2X1 i_1454 ( .Y (n_1618),
	.B (n_911),
	.A (n_2382) );
   AOI211X1 i_361 ( .Y (n_1617),
	.C0 (n_1616),
	.B0 (n_1827),
	.A1 (n_1831),
	.A0 (n_1830) );
   NOR2X1 i_1451 ( .Y (n_1616),
	.B (n_1880),
	.A (n_906) );
   NOR2X1 i_1449 ( .Y (n_1614),
	.B (op_a[27]),
	.A (n_1936) );
   NAND2BX1 i_1448 ( .Y (n_1613),
	.B (n_3062),
	.AN (n_949) );
   NAND3X1 i_446 ( .Y (n_1612),
	.C (n_1754),
	.B (n_1611),
	.A (n_879) );
   NAND3BX1 i_1445 ( .Y (n_1611),
	.C (n_946),
	.B (n_1758),
	.AN (n_1806) );
   OAI21XL i_778553 ( .Y (result[26]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1609) );
   AOI211X1 i_1351 ( .Y (n_1609),
	.C0 (n_2378),
	.B0 (n_1727),
	.A1 (n_2360),
	.A0 (n_1598) );
   OAI21XL i_261 ( .Y (n_1600),
	.B0 (n_1596),
	.A1 (n_1699),
	.A0 (n_2370) );
   AOI21X1 i_262 ( .Y (n_1599),
	.B0 (n_1589),
	.A1 (n_2372),
	.A0 (op_a[26]) );
   OAI2BB1X1 i_263 ( .Y (n_1598),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1708) );
   NAND2X1 i_1424 ( .Y (n_1596),
	.B (n_2370),
	.A (n_1699) );
   AOI211X1 i_356 ( .Y (n_1594),
	.C0 (n_1593),
	.B0 (n_2299),
	.A1 (n_2300),
	.A0 (n_2264) );
   NOR4BX1 i_1419 ( .Y (n_1593),
	.D (n_1494),
	.C (n_1395),
	.B (n_1441),
	.AN (n_2300) );
   NOR2X1 i_251379 ( .Y (n_1592),
	.B (op_a[25]),
	.A (op_b[25]) );
   NOR2X1 i_1416 ( .Y (n_1589),
	.B (op_a[26]),
	.A (n_2372) );
   OAI211X1 i_445 ( .Y (n_1587),
	.C0 (n_1586),
	.B0 (n_2294),
	.A1 (n_2259),
	.A0 (n_2295) );
   NAND4BXL i_1410 ( .Y (n_1586),
	.D (n_1487),
	.C (n_925),
	.B (n_1485),
	.AN (n_2260) );
   NAND2BX1 i_577104 ( .Y (n_1585),
	.B (op_b[25]),
	.AN (op_a[25]) );
   OAI21XL i_788554 ( .Y (result[25]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1582) );
   AOI211X1 i_1342 ( .Y (n_1582),
	.C0 (n_2358),
	.B0 (n_1727),
	.A1 (n_2341),
	.A0 (n_1571) );
   NOR2X1 i_1384 ( .Y (n_1579),
	.B (n_3095),
	.A (n_1573) );
   AOI31X1 i_252 ( .Y (n_1573),
	.B0 (n_1568),
	.A2 (n_2349),
	.A1 (n_2346),
	.A0 (n_1566) );
   AOI31X1 i_253 ( .Y (n_1572),
	.B0 (n_1563),
	.A2 (n_2351),
	.A1 (op_a[25]),
	.A0 (n_2285) );
   OAI21XL i_254 ( .Y (n_1571),
	.B0 (n_1716),
	.A1 (n_1738),
	.A0 (n_2344) );
   AOI21X1 i_1375 ( .Y (n_1568),
	.B0 (n_2349),
	.A1 (n_2346),
	.A0 (n_1566) );
   AOI211X1 i_355 ( .Y (n_1567),
	.C0 (n_1565),
	.B0 (n_1830),
	.A1 (n_1879),
	.A0 (n_1835) );
   NAND3BX1 i_1373 ( .Y (n_1566),
	.C (n_1831),
	.B (n_1881),
	.AN (n_1567) );
   NOR4BX1 i_1371 ( .Y (n_1565),
	.D (n_1467),
	.C (n_1390),
	.B (n_1395),
	.AN (n_1879) );
   AOI21X1 i_1368 ( .Y (n_1563),
	.B0 (op_a[25]),
	.A1 (n_2285),
	.A0 (n_2351) );
   OAI211X1 i_444 ( .Y (n_1561),
	.C0 (n_1559),
	.B0 (n_1757),
	.A1 (n_1762),
	.A0 (n_1806) );
   NAND4BXL i_1361 ( .Y (n_1559),
	.D (n_1383),
	.C (n_927),
	.B (n_1462),
	.AN (n_1806) );
   OAI21XL i_798555 ( .Y (result[24]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1557) );
   AOI211X1 i_1333 ( .Y (n_1557),
	.C0 (n_2339),
	.B0 (n_1727),
	.A1 (n_2323),
	.A0 (n_1546) );
   OAI21XL i_245 ( .Y (n_1548),
	.B0 (n_1543),
	.A1 (n_1647),
	.A0 (n_2333) );
   AOI21X1 i_246 ( .Y (n_1547),
	.B0 (n_1536),
	.A1 (n_1907),
	.A0 (op_a[24]) );
   OAI2BB1X1 i_248 ( .Y (n_1546),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1637) );
   NOR2X1 i_241378 ( .Y (n_1544),
	.B (op_a[24]),
	.A (op_b[24]) );
   NAND2X1 i_1338 ( .Y (n_1543),
	.B (n_2333),
	.A (n_1647) );
   AOI211X1 i_354 ( .Y (n_1541),
	.C0 (n_1540),
	.B0 (n_2264),
	.A1 (n_2265),
	.A0 (n_2233) );
   NOR4BX1 i_1332 ( .Y (n_1540),
	.D (n_1443),
	.C (n_1395),
	.B (n_1441),
	.AN (n_2234) );
   NOR2X1 i_231377 ( .Y (n_1539),
	.B (op_a[23]),
	.A (op_b[23]) );
   NOR2X1 i_1329 ( .Y (n_1536),
	.B (op_a[24]),
	.A (n_1907) );
   OAI211X1 i_437 ( .Y (n_1534),
	.C0 (n_1533),
	.B0 (n_2259),
	.A1 (n_2260),
	.A0 (n_2228) );
   NAND4BXL i_1323 ( .Y (n_1533),
	.D (n_929),
	.C (n_1436),
	.B (n_1383),
	.AN (n_2260) );
   NAND2BX1 i_557102 ( .Y (n_1532),
	.B (op_b[23]),
	.AN (op_a[23]) );
   OAI21XL i_808556 ( .Y (result[23]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1529) );
   AOI211X1 i_1324 ( .Y (n_1529),
	.C0 (n_2321),
	.B0 (n_1727),
	.A1 (n_2313),
	.A0 (n_1518) );
   OAI21XL i_238 ( .Y (n_1520),
	.B0 (n_1516),
	.A1 (n_1617),
	.A0 (n_2315) );
   AOI31X1 i_240 ( .Y (n_1519),
	.B0 (n_1513),
	.A2 (n_1932),
	.A1 (op_a[23]),
	.A0 (n_1930) );
   OAI2BB1X1 i_241 ( .Y (n_1518),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1612) );
   NAND2X1 i_1300 ( .Y (n_1516),
	.B (n_2315),
	.A (n_1617) );
   AOI21X1 i_1296 ( .Y (n_1513),
	.B0 (op_a[23]),
	.A1 (n_1930),
	.A0 (n_1932) );
   OAI21XL i_818557 ( .Y (result[22]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1510) );
   AOI211X1 i_1315 ( .Y (n_1510),
	.C0 (n_2311),
	.B0 (n_1727),
	.A1 (n_2293),
	.A0 (n_1499) );
   OAI21XL i_232 ( .Y (n_1501),
	.B0 (n_1496),
	.A1 (n_1594),
	.A0 (n_2303) );
   XNOR2X1 i_233 ( .Y (n_1500),
	.B (n_2305),
	.A (op_a[22]) );
   OAI2BB1X1 i_234 ( .Y (n_1499),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1587) );
   NOR2X1 i_221376 ( .Y (n_1497),
	.B (op_a[22]),
	.A (op_b[22]) );
   NAND2X1 i_1273 ( .Y (n_1496),
	.B (n_2303),
	.A (n_1594) );
   AOI211X1 i_352 ( .Y (n_1494),
	.C0 (n_1493),
	.B0 (n_2233),
	.A1 (n_2234),
	.A0 (n_2198) );
   NOR4BX1 i_1267 ( .Y (n_1493),
	.D (n_1392),
	.C (n_1297),
	.B (n_1339),
	.AN (n_2234) );
   NOR2X1 i_211375 ( .Y (n_1492),
	.B (op_a[21]),
	.A (op_b[21]) );
   OAI211X1 i_435 ( .Y (n_1487),
	.C0 (n_1486),
	.B0 (n_2228),
	.A1 (n_2193),
	.A0 (n_2229) );
   NAND4BXL i_1257 ( .Y (n_1486),
	.D (n_1385),
	.C (n_929),
	.B (n_1383),
	.AN (n_2194) );
   NAND2BX1 i_537100 ( .Y (n_1485),
	.B (op_b[21]),
	.AN (op_a[21]) );
   OAI21XL i_828558 ( .Y (result[21]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1482) );
   AOI211X1 i_1306 ( .Y (n_1482),
	.C0 (n_2291),
	.B0 (n_1727),
	.A1 (n_2276),
	.A0 (n_1471) );
   OAI21XL i_225 ( .Y (n_1473),
	.B0 (n_1469),
	.A1 (n_1567),
	.A0 (n_2282) );
   AOI21X1 i_226 ( .Y (n_1472),
	.B0 (n_1464),
	.A1 (n_2285),
	.A0 (op_a[21]) );
   OAI2BB1X1 i_228 ( .Y (n_1471),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1561) );
   NAND2X1 i_1233 ( .Y (n_1469),
	.B (n_2282),
	.A (n_1567) );
   AOI211X1 i_351 ( .Y (n_1467),
	.C0 (n_1466),
	.B0 (n_1838),
	.A1 (n_1877),
	.A0 (n_1843) );
   NOR4BX1 i_1228 ( .Y (n_1466),
	.D (n_1365),
	.C (n_1293),
	.B (n_1297),
	.AN (n_1877) );
   NOR2X1 i_1226 ( .Y (n_1464),
	.B (op_a[21]),
	.A (n_2285) );
   OAI211X1 i_434 ( .Y (n_1462),
	.C0 (n_1461),
	.B0 (n_1765),
	.A1 (n_1770),
	.A0 (n_1804) );
   NAND4BXL i_1218 ( .Y (n_1461),
	.D (n_1286),
	.C (n_931),
	.B (n_1360),
	.AN (n_1804) );
   OAI21XL i_838559 ( .Y (result[20]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1459) );
   AOI211X1 i_1297 ( .Y (n_1459),
	.C0 (n_2274),
	.B0 (n_1727),
	.A1 (n_2258),
	.A0 (n_1448) );
   OAI21XL i_217 ( .Y (n_1450),
	.B0 (n_1445),
	.A1 (n_1541),
	.A0 (n_2268) );
   XNOR2X1 i_218 ( .Y (n_1449),
	.B (n_1903),
	.A (op_a[20]) );
   OAI2BB1X1 i_219 ( .Y (n_1448),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1534) );
   NOR2X1 i_201374 ( .Y (n_1446),
	.B (op_a[20]),
	.A (op_b[20]) );
   NAND2X1 i_1195 ( .Y (n_1445),
	.B (n_2268),
	.A (n_1541) );
   AOI211X1 i_350 ( .Y (n_1443),
	.C0 (n_1442),
	.B0 (n_2198),
	.A1 (n_2199),
	.A0 (n_2167) );
   NOR4BX1 i_1190 ( .Y (n_1442),
	.D (n_1340),
	.C (n_1297),
	.B (n_1339),
	.AN (n_2168) );
   NOR2X1 i_191373 ( .Y (n_1441),
	.B (op_a[19]),
	.A (op_b[19]) );
   OAI211X1 i_433 ( .Y (n_1436),
	.C0 (n_1435),
	.B0 (n_2193),
	.A1 (n_2194),
	.A0 (n_2162) );
   NAND4BXL i_1181 ( .Y (n_1435),
	.D (n_933),
	.C (n_1334),
	.B (n_1286),
	.AN (n_2194) );
   NAND2BX1 i_517098 ( .Y (n_1434),
	.B (op_b[19]),
	.AN (op_a[19]) );
   OAI21XL i_848560 ( .Y (result[19]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1431) );
   AOI211X1 i_1288 ( .Y (n_1431),
	.C0 (n_2256),
	.B0 (n_1727),
	.A1 (n_2248),
	.A0 (n_1420) );
   OAI21XL i_167 ( .Y (n_1422),
	.B0 (n_1418),
	.A1 (n_906),
	.A0 (n_2250) );
   AOI21X1 i_186 ( .Y (n_1421),
	.B0 (n_1413),
	.A1 (n_1930),
	.A0 (op_a[19]) );
   OAI2BB1X1 i_188 ( .Y (n_1420),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_946) );
   NAND2X1 i_1157 ( .Y (n_1418),
	.B (n_2250),
	.A (n_906) );
   AOI211X1 i_348 ( .Y (n_1416),
	.C0 (n_1415),
	.B0 (n_1843),
	.A1 (n_1847),
	.A0 (n_1846) );
   NOR4BX1 i_1151 ( .Y (n_1415),
	.D (n_903),
	.C (n_1293),
	.B (n_1297),
	.AN (n_1875) );
   NOR2X1 i_1149 ( .Y (n_1413),
	.B (op_a[19]),
	.A (n_1930) );
   OAI211X1 i_432 ( .Y (n_1411),
	.C0 (n_1410),
	.B0 (n_1770),
	.A1 (n_1774),
	.A0 (n_1773) );
   NAND4BXL i_1143 ( .Y (n_1410),
	.D (n_943),
	.C (n_1286),
	.B (n_931),
	.AN (n_1802) );
   OAI21XL i_858561 ( .Y (result[18]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1408) );
   AOI211X1 i_1279 ( .Y (n_1408),
	.C0 (n_2246),
	.B0 (n_1727),
	.A1 (n_2227),
	.A0 (n_1397) );
   OAI21XL i_130 ( .Y (n_1399),
	.B0 (n_1394),
	.A1 (n_1494),
	.A0 (n_2237) );
   AOI31X1 i_131 ( .Y (n_1398),
	.B0 (n_1387),
	.A2 (n_2239),
	.A1 (op_a[18]),
	.A0 (n_2174) );
   OAI2BB1X1 i_132 ( .Y (n_1397),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1487) );
   NOR2X1 i_181372 ( .Y (n_1395),
	.B (op_a[18]),
	.A (op_b[18]) );
   NAND2X1 i_1121 ( .Y (n_1394),
	.B (n_2237),
	.A (n_1494) );
   AOI211X1 i_347 ( .Y (n_1392),
	.C0 (n_1391),
	.B0 (n_2167),
	.A1 (n_2168),
	.A0 (n_2132) );
   NOR4BX1 i_1115 ( .Y (n_1391),
	.D (n_1294),
	.C (n_1198),
	.B (n_1244),
	.AN (n_2168) );
   NOR2X1 i_171371 ( .Y (n_1390),
	.B (op_a[17]),
	.A (op_b[17]) );
   AOI21X1 i_1112 ( .Y (n_1387),
	.B0 (op_a[18]),
	.A1 (n_2174),
	.A0 (n_2239) );
   OAI211X1 i_431 ( .Y (n_1385),
	.C0 (n_1384),
	.B0 (n_2162),
	.A1 (n_2127),
	.A0 (n_2163) );
   NAND4BXL i_1105 ( .Y (n_1384),
	.D (n_1287),
	.C (n_933),
	.B (n_1286),
	.AN (n_2128) );
   NAND2BX1 i_497096 ( .Y (n_1383),
	.B (op_b[17]),
	.AN (op_a[17]) );
   OAI21XL i_868562 ( .Y (result[17]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1380) );
   AOI211X1 i_1270 ( .Y (n_1380),
	.C0 (n_2225),
	.B0 (n_1727),
	.A1 (n_2210),
	.A0 (n_1369) );
   OAI21XL i_125 ( .Y (n_1371),
	.B0 (n_1367),
	.A1 (n_1467),
	.A0 (n_2216) );
   AOI31X1 i_126 ( .Y (n_1370),
	.B0 (n_1362),
	.A2 (n_2218),
	.A1 (op_a[17]),
	.A0 (n_2153) );
   OAI2BB1X1 i_127 ( .Y (n_1369),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1462) );
   NAND2X1 i_1075 ( .Y (n_1367),
	.B (n_2216),
	.A (n_1467) );
   AOI211X1 i_346 ( .Y (n_1365),
	.C0 (n_1364),
	.B0 (n_1846),
	.A1 (n_1875),
	.A0 (n_1851) );
   NOR4BX1 i_1070 ( .Y (n_1364),
	.D (n_1268),
	.C (n_1193),
	.B (n_1198),
	.AN (n_1875) );
   AOI21X1 i_1068 ( .Y (n_1362),
	.B0 (op_a[17]),
	.A1 (n_2153),
	.A0 (n_2218) );
   OAI211X1 i_430 ( .Y (n_1360),
	.C0 (n_1359),
	.B0 (n_1773),
	.A1 (n_1778),
	.A0 (n_1802) );
   NAND4BXL i_1061 ( .Y (n_1359),
	.D (n_1186),
	.C (n_935),
	.B (n_1264),
	.AN (n_1802) );
   OAI21XL i_878563 ( .Y (result[16]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1357) );
   AOI211X1 i_1261 ( .Y (n_1357),
	.C0 (n_2208),
	.B0 (n_1727),
	.A1 (n_2192),
	.A0 (n_1346) );
   OAI21XL i_120 ( .Y (n_1348),
	.B0 (n_1343),
	.A1 (n_1443),
	.A0 (n_2202) );
   AOI21X1 i_121 ( .Y (n_1347),
	.B0 (n_1337),
	.A1 (n_1899),
	.A0 (op_a[16]) );
   OAI2BB1X1 i_122 ( .Y (n_1346),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1436) );
   NOR2X1 i_161370 ( .Y (n_1344),
	.B (op_a[16]),
	.A (op_b[16]) );
   NAND2X1 i_1041 ( .Y (n_1343),
	.B (n_2202),
	.A (n_1443) );
   NOR4BX1 i_345 ( .Y (n_1341),
	.D (n_1245),
	.C (n_1198),
	.B (n_1244),
	.AN (n_2103) );
   AOI211X1 i_1038 ( .Y (n_1340),
	.C0 (n_1341),
	.B0 (n_2132),
	.A1 (n_2133),
	.A0 (n_2102) );
   NOR2X1 i_151369 ( .Y (n_1339),
	.B (op_a[15]),
	.A (op_b[15]) );
   NOR2X1 i_1035 ( .Y (n_1337),
	.B (op_a[16]),
	.A (n_1899) );
   OAI211X1 i_429 ( .Y (n_1334),
	.C0 (n_1333),
	.B0 (n_2127),
	.A1 (n_2128),
	.A0 (n_2097) );
   NAND4BXL i_1029 ( .Y (n_1333),
	.D (n_937),
	.C (n_1238),
	.B (n_1186),
	.AN (n_2128) );
   NAND2BX1 i_477094 ( .Y (n_1332),
	.B (op_b[15]),
	.AN (op_a[15]) );
   OAI21XL i_888564 ( .Y (result[15]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1329) );
   AOI211X1 i_1252 ( .Y (n_1329),
	.C0 (n_2190),
	.B0 (n_1727),
	.A1 (n_2182),
	.A0 (n_1318) );
   OAI21XL i_115 ( .Y (n_1320),
	.B0 (n_1316),
	.A1 (n_1416),
	.A0 (n_2184) );
   AOI31X1 i_116 ( .Y (n_1319),
	.B0 (n_1314),
	.A2 (n_1926),
	.A1 (op_a[15]),
	.A0 (n_1924) );
   OAI2BB1X1 i_117 ( .Y (n_1318),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1411) );
   NAND2X1 i_1008 ( .Y (n_1316),
	.B (n_2184),
	.A (n_1416) );
   AOI21X1 i_1006 ( .Y (n_1314),
	.B0 (op_a[15]),
	.A1 (n_1924),
	.A0 (n_1926) );
   OAI21XL i_898565 ( .Y (result[14]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1310) );
   AOI211X1 i_1243 ( .Y (n_1310),
	.C0 (n_2180),
	.B0 (n_1727),
	.A1 (n_2161),
	.A0 (n_1299) );
   OAI21XL i_110 ( .Y (n_1301),
	.B0 (n_1296),
	.A1 (n_1392),
	.A0 (n_2171) );
   AOI21X1 i_111 ( .Y (n_1300),
	.B0 (n_1291),
	.A1 (n_2174),
	.A0 (op_a[14]) );
   OAI2BB1X1 i_112 ( .Y (n_1299),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1385) );
   NOR2X1 i_141368 ( .Y (n_1297),
	.B (op_a[14]),
	.A (op_b[14]) );
   NAND2X1 i_984 ( .Y (n_1296),
	.B (n_2171),
	.A (n_1392) );
   AOI211X1 i_981 ( .Y (n_1294),
	.C0 (n_855),
	.B0 (n_2102),
	.A1 (n_2103),
	.A0 (n_2066) );
   NOR2X1 i_131367 ( .Y (n_1293),
	.B (op_a[13]),
	.A (op_b[13]) );
   NOR2X1 i_978 ( .Y (n_1291),
	.B (op_a[14]),
	.A (n_2174) );
   NAND4X1 i_426 ( .Y (n_1288),
	.D (n_2062),
	.C (n_1187),
	.B (n_937),
	.A (n_1186) );
   OAI211X1 i_972 ( .Y (n_1287),
	.C0 (n_1288),
	.B0 (n_2097),
	.A1 (n_2061),
	.A0 (n_2098) );
   NAND2BX1 i_457092 ( .Y (n_1286),
	.B (op_b[13]),
	.AN (op_a[13]) );
   OAI21XL i_908566 ( .Y (result[13]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1283) );
   AOI211X1 i_1234 ( .Y (n_1283),
	.C0 (n_2159),
	.B0 (n_1727),
	.A1 (n_2144),
	.A0 (n_1272) );
   OAI21XL i_105 ( .Y (n_1274),
	.B0 (n_1270),
	.A1 (n_1365),
	.A0 (n_2150) );
   AOI21X1 i_106 ( .Y (n_1273),
	.B0 (n_1267),
	.A1 (n_2153),
	.A0 (op_a[13]) );
   OAI2BB1X1 i_107 ( .Y (n_1272),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1360) );
   NAND2X1 i_950 ( .Y (n_1270),
	.B (n_2150),
	.A (n_1365) );
   AOI31X1 i_947 ( .Y (n_1268),
	.B0 (n_3092),
	.A2 (n_1167),
	.A1 (n_1863),
	.A0 (n_1873) );
   NOR2X1 i_945 ( .Y (n_1267),
	.B (op_a[13]),
	.A (n_2153) );
   OAI31X1 i_939 ( .Y (n_1264),
	.B0 (n_2080),
	.A2 (n_1162),
	.A1 (n_1790),
	.A0 (n_1800) );
   OAI21XL i_918567 ( .Y (result[12]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1262) );
   AOI211X1 i_1225 ( .Y (n_1262),
	.C0 (n_2142),
	.B0 (n_1727),
	.A1 (n_2126),
	.A0 (n_1251) );
   OAI21XL i_99 ( .Y (n_1253),
	.B0 (n_1248),
	.A1 (n_1340),
	.A0 (n_2136) );
   XNOR2X1 i_100 ( .Y (n_1252),
	.B (op_a[12]),
	.A (n_1895) );
   OAI2BB1X1 i_101 ( .Y (n_1251),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1334) );
   NOR2X1 i_121366 ( .Y (n_1249),
	.B (op_a[12]),
	.A (op_b[12]) );
   NAND2X1 i_918 ( .Y (n_1248),
	.B (n_2136),
	.A (n_1340) );
   NOR4BX1 i_336 ( .Y (n_1246),
	.D (n_2004),
	.C (n_1100),
	.B (n_1144),
	.AN (n_2039) );
   AOI211X1 i_915 ( .Y (n_1245),
	.C0 (n_1246),
	.B0 (n_2066),
	.A1 (n_2067),
	.A0 (n_2038) );
   NOR2X1 i_111365 ( .Y (n_1244),
	.B (op_a[11]),
	.A (op_b[11]) );
   NAND4X1 i_422 ( .Y (n_1239),
	.D (n_942),
	.C (n_1137),
	.B (n_2062),
	.A (n_1090) );
   NAND3X1 i_908 ( .Y (n_1238),
	.C (n_862),
	.B (n_1239),
	.A (n_2061) );
   NAND2BX1 i_437090 ( .Y (n_1237),
	.B (op_b[11]),
	.AN (op_a[11]) );
   OAI21XL i_928568 ( .Y (result[11]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1234) );
   AOI211X1 i_1216 ( .Y (n_1234),
	.C0 (n_2124),
	.B0 (n_1727),
	.A1 (n_2116),
	.A0 (n_1223) );
   OAI21XL i_94 ( .Y (n_1225),
	.B0 (n_1221),
	.A1 (n_903),
	.A0 (n_2118) );
   AOI21X1 i_95 ( .Y (n_1224),
	.B0 (n_1217),
	.A1 (n_1924),
	.A0 (op_a[11]) );
   OAI2BB1X1 i_96 ( .Y (n_1223),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_943) );
   NAND2X1 i_886 ( .Y (n_1221),
	.B (n_2118),
	.A (n_903) );
   NOR4BX1 i_334 ( .Y (n_1219),
	.D (n_1870),
	.C (n_1097),
	.B (n_1053),
	.AN (n_1863) );
   AOI211X1 i_883 ( .Y (n_1218),
	.C0 (n_1219),
	.B0 (n_1859),
	.A1 (n_1863),
	.A0 (n_1862) );
   NOR2X1 i_881 ( .Y (n_1217),
	.B (op_a[11]),
	.A (n_1924) );
   AOI211X1 i_877 ( .Y (n_1213),
	.C0 (n_1786),
	.B0 (n_861),
	.A1 (n_1799),
	.A0 (n_1797) );
   OAI21XL i_938569 ( .Y (result[10]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1211) );
   AOI211X1 i_1207 ( .Y (n_1211),
	.C0 (n_2114),
	.B0 (n_1727),
	.A1 (n_2096),
	.A0 (n_1200) );
   OAI21XL i_89 ( .Y (n_1202),
	.B0 (n_1197),
	.A1 (n_1294),
	.A0 (n_2106) );
   AOI21X1 i_90 ( .Y (n_1201),
	.B0 (n_1191),
	.A1 (n_2108),
	.A0 (op_a[10]) );
   OAI2BB1X1 i_91 ( .Y (n_1200),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1287) );
   NOR2X1 i_101364 ( .Y (n_1198),
	.B (op_a[10]),
	.A (op_b[10]) );
   NAND2X1 i_856 ( .Y (n_1197),
	.B (n_2106),
	.A (n_1294) );
   AOI31X1 i_853 ( .Y (n_1194),
	.B0 (n_3089),
	.A2 (n_1976),
	.A1 (n_2003),
	.A0 (n_2039) );
   NOR2X1 i_91363 ( .Y (n_1193),
	.B (op_a[9]),
	.A (op_b[9]) );
   NOR2X1 i_851 ( .Y (n_1191),
	.B (op_a[10]),
	.A (n_2108) );
   NAND4BXL i_418 ( .Y (n_1188),
	.D (n_1972),
	.C (n_942),
	.B (n_1090),
	.AN (n_1997) );
   NAND4X1 i_846 ( .Y (n_1187),
	.D (n_860),
	.C (n_1188),
	.B (n_1785),
	.A (n_1089) );
   NAND2BX1 i_417088 ( .Y (n_1186),
	.B (op_b[9]),
	.AN (op_a[9]) );
   OAI21XL i_948570 ( .Y (result[9]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1183) );
   AOI211X1 i_1198 ( .Y (n_1183),
	.C0 (n_2094),
	.B0 (n_1727),
	.A1 (n_2079),
	.A0 (n_1172) );
   OAI21XL i_84 ( .Y (n_1174),
	.B0 (n_1170),
	.A1 (n_1268),
	.A0 (n_2085) );
   AOI31X1 i_85 ( .Y (n_1173),
	.B0 (n_1166),
	.A2 (n_2087),
	.A1 (op_a[9]),
	.A0 (n_2017) );
   OAI2BB1X1 i_86 ( .Y (n_1172),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1264) );
   NAND2X1 i_824 ( .Y (n_1170),
	.B (n_2085),
	.A (n_1268) );
   NAND3X1 i_18 ( .Y (n_1168),
	.C (n_1871),
	.B (n_3085),
	.A (n_1869) );
   NAND2X1 i_821 ( .Y (n_1167),
	.B (n_2020),
	.A (n_1168) );
   AOI21X1 i_820 ( .Y (n_1166),
	.B0 (op_a[9]),
	.A1 (n_2017),
	.A0 (n_2087) );
   AOI2BB1X1 i_814 ( .Y (n_1162),
	.B0 (n_2013),
	.A1N (n_857),
	.A0N (n_1798) );
   OAI21XL i_958571 ( .Y (result[8]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1160) );
   AOI211X1 i_1189 ( .Y (n_1160),
	.C0 (n_2077),
	.B0 (n_1727),
	.A1 (n_2060),
	.A0 (n_1149) );
   OAI21XL i_79 ( .Y (n_1151),
	.B0 (n_1146),
	.A1 (n_1245),
	.A0 (n_2070) );
   XNOR2X1 i_80 ( .Y (n_1150),
	.B (n_1891),
	.A (op_a[8]) );
   OAI2BB1X1 i_81 ( .Y (n_1149),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1238) );
   NOR2X1 i_81362 ( .Y (n_1147),
	.B (op_a[8]),
	.A (op_b[8]) );
   NAND2X1 i_794 ( .Y (n_1146),
	.B (n_2070),
	.A (n_1245) );
   NOR2X1 i_7 ( .Y (n_1144),
	.B (op_a[7]),
	.A (op_b[7]) );
   OAI21XL i_784 ( .Y (n_1137),
	.B0 (n_1998),
	.A1 (n_1997),
	.A0 (n_856) );
   NOR2BX1 i_337080 ( .Y (n_1136),
	.B (op_a[1]),
	.AN (op_b[1]) );
   NAND2BX1 i_397086 ( .Y (n_1135),
	.B (op_b[7]),
	.AN (op_a[7]) );
   OAI21XL i_968572 ( .Y (result[7]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1132) );
   AOI21X1 i_1180 ( .Y (n_1132),
	.B0 (n_2059),
	.A1 (n_2049),
	.A0 (n_1122) );
   AOI21X1 i_768 ( .Y (n_1129),
	.B0 (n_1917),
	.A1 (n_2052),
	.A0 (n_1915) );
   OAI21XL i_73 ( .Y (n_1123),
	.B0 (n_1119),
	.A1 (n_1218),
	.A0 (n_2053) );
   OAI2BB1X1 i_74 ( .Y (n_1122),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_3076) );
   NAND2X1 i_763 ( .Y (n_1119),
	.B (n_2053),
	.A (n_1218) );
   NOR2X1 i_759 ( .Y (n_1116),
	.B (n_2051),
	.A (op_a[7]) );
   OAI21XL i_978573 ( .Y (result[6]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1113) );
   AOI21X1 i_1171 ( .Y (n_1113),
	.B0 (n_2048),
	.A1 (n_2028),
	.A0 (n_1103) );
   AOI21X1 i_744 ( .Y (n_1110),
	.B0 (n_1917),
	.A1 (n_2037),
	.A0 (n_1915) );
   OAI21XL i_66 ( .Y (n_1104),
	.B0 (n_1099),
	.A1 (n_1194),
	.A0 (n_2042) );
   OAI2BB1X1 i_67 ( .Y (n_1103),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1187) );
   NOR2X1 i_61361 ( .Y (n_1100),
	.B (op_a[6]),
	.A (op_b[6]) );
   NAND2X1 i_739 ( .Y (n_1099),
	.B (n_2042),
	.A (n_1194) );
   NOR2X1 i_31360 ( .Y (n_1097),
	.B (op_a[3]),
	.A (op_b[3]) );
   NOR2X1 i_21359 ( .Y (n_1096),
	.B (op_a[2]),
	.A (op_b[2]) );
   NOR2X1 i_5 ( .Y (n_1095),
	.B (op_a[5]),
	.A (op_b[5]) );
   NOR2X1 i_732 ( .Y (n_1092),
	.B (n_2036),
	.A (op_a[6]) );
   NAND2BX1 i_377084 ( .Y (n_1090),
	.B (op_b[5]),
	.AN (op_a[5]) );
   NAND2X1 i_726 ( .Y (n_1089),
	.B (n_1787),
	.A (n_1090) );
   OAI21XL i_988574 ( .Y (result[5]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1087) );
   NOR4BX1 i_1162 ( .Y (n_1087),
	.D (n_1076),
	.C (n_2025),
	.B (n_1084),
	.AN (n_1085) );
   NAND4X1 i_715 ( .Y (n_1085),
	.D (n_3062),
	.C (n_1162),
	.B (n_1090),
	.A (n_1785) );
   AOI21X1 i_712 ( .Y (n_1084),
	.B0 (n_1917),
	.A1 (n_2019),
	.A0 (n_1915) );
   AOI31X1 i_60 ( .Y (n_1078),
	.B0 (n_1073),
	.A2 (n_2021),
	.A1 (n_2020),
	.A0 (n_1168) );
   AOI22X1 i_713 ( .Y (n_1076),
	.B1 (n_1090),
	.B0 (n_1785),
	.A1 (n_1071),
	.A0 (n_1716) );
   AOI21X1 i_706 ( .Y (n_1073),
	.B0 (n_2021),
	.A1 (n_2020),
	.A0 (n_1168) );
   NOR2X1 i_1 ( .Y (n_1072),
	.B (op_a[1]),
	.A (op_b[1]) );
   NAND2BX1 i_703 ( .Y (n_1071),
	.B (n_3062),
	.AN (n_1162) );
   NOR2X1 i_701 ( .Y (n_1070),
	.B (n_2018),
	.A (op_a[5]) );
   NAND2BX1 i_347081 ( .Y (n_1068),
	.B (op_b[2]),
	.AN (op_a[2]) );
   OAI21XL i_998575 ( .Y (result[4]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1066) );
   AOI21X1 i_1153 ( .Y (n_1066),
	.B0 (n_2011),
	.A1 (n_1995),
	.A0 (n_1056) );
   AOI21X1 i_681 ( .Y (n_1063),
	.B0 (n_1917),
	.A1 (n_2001),
	.A0 (n_1915) );
   OAI21XL i_55 ( .Y (n_1057),
	.B0 (n_1052),
	.A1 (n_2004),
	.A0 (n_2005) );
   OAI2BB1X1 i_56 ( .Y (n_1056),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1137) );
   NOR2X1 i_4 ( .Y (n_1053),
	.B (op_a[4]),
	.A (op_b[4]) );
   NAND2X1 i_676 ( .Y (n_1052),
	.B (n_2005),
	.A (n_2004) );
   NOR2X1 i_670 ( .Y (n_1048),
	.B (n_2000),
	.A (op_a[4]) );
   NAND2BX1 i_357082 ( .Y (n_1045),
	.B (op_b[3]),
	.AN (op_a[3]) );
   OAI21XL i_1008576 ( .Y (result[3]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1042) );
   AOI21X1 i_1144 ( .Y (n_1042),
	.B0 (n_1994),
	.A1 (n_1984),
	.A0 (n_1032) );
   AOI21X1 i_651 ( .Y (n_1039),
	.B0 (n_1917),
	.A1 (n_1987),
	.A0 (n_1915) );
   OAI21XL i_49 ( .Y (n_1033),
	.B0 (n_1029),
	.A1 (n_1870),
	.A0 (n_1988) );
   OAI2BB1X1 i_50 ( .Y (n_1032),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1797) );
   NAND2X1 i_646 ( .Y (n_1029),
	.B (n_1988),
	.A (n_1870) );
   NOR2X1 i_642 ( .Y (n_1026),
	.B (n_1986),
	.A (op_a[3]) );
   OAI21XL i_1018577 ( .Y (result[2]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1023) );
   AOI21X1 i_1135 ( .Y (n_1023),
	.B0 (n_1983),
	.A1 (n_1970),
	.A0 (n_1013) );
   AOI21X1 i_627 ( .Y (n_1020),
	.B0 (n_1917),
	.A1 (n_1975),
	.A0 (n_1915) );
   XOR2X1 i_43 ( .Y (n_1014),
	.B (n_1977),
	.A (n_1976) );
   OAI2BB1X1 i_44 ( .Y (n_1013),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1972) );
   NOR2X1 i_617 ( .Y (n_1006),
	.B (n_1974),
	.A (op_a[2]) );
   OAI21XL i_1028578 ( .Y (result[1]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1002) );
   AOI21X1 i_1126 ( .Y (n_1002),
	.B0 (n_1969),
	.A1 (n_1959),
	.A0 (n_992) );
   AOI21X1 i_601 ( .Y (n_999),
	.B0 (n_1917),
	.A1 (n_1962),
	.A0 (n_1915) );
   OAI31X1 i_37 ( .Y (n_993),
	.B0 (n_988),
	.A2 (n_3085),
	.A1 (n_1072),
	.A0 (n_3083) );
   OAI2BB1X1 i_38 ( .Y (n_992),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_1795) );
   OAI21XL i_595 ( .Y (n_988),
	.B0 (n_3085),
	.A1 (n_3083),
	.A0 (n_1072) );
   NOR2X1 i_592 ( .Y (n_986),
	.B (n_1961),
	.A (op_a[1]) );
   AOI21X1 i_1038579 ( .Y (n_984),
	.B0 (n_827),
	.A1 (n_9076575),
	.A0 (n_983) );
   NAND3BX1 i_1117 ( .Y (n_983),
	.C (n_976),
	.B (n_1957),
	.AN (n_981) );
   AOI21X1 i_582 ( .Y (n_981),
	.B0 (n_1795),
	.A1 (n_1738),
	.A0 (n_1716) );
   OR2X1 i_34 ( .Y (n_978),
	.B (n_974),
	.A (n_1946) );
   OAI21XL i_583 ( .Y (n_976),
	.B0 (op_a[0]),
	.A1 (n_1955),
	.A0 (n_973) );
   NOR2X1 i_574 ( .Y (n_974),
	.B (n_3095),
	.A (n_3085) );
   AOI21X1 i_575 ( .Y (n_973),
	.B0 (op_b[0]),
	.A1 (n_1738),
	.A0 (n_1716) );
   NOR3X1 i_570 ( .Y (n_971),
	.C (n_1733),
	.B (op_a[31]),
	.A (n_1950) );
   NOR2X1 i_569 ( .Y (n_970),
	.B (n_3095),
	.A (op_b[31]) );
   NAND4X1 i_559 ( .Y (n_967),
	.D (n_1918),
	.C (n_1938),
	.B (n_1915),
	.A (n_1936) );
   AOI22X1 i_291 ( .Y (n_964),
	.B1 (n_868),
	.B0 (n_1883),
	.A1 (n_3062),
	.A0 (n_1810) );
   NAND3X1 i_292 ( .Y (n_963),
	.C (n_1942),
	.B (n_1944),
	.A (n_958) );
   OAI221XL i_293 ( .Y (n_962),
	.C0 (n_1716),
	.B1 (n_1738),
	.B0 (n_1810),
	.A1 (n_1883),
	.A0 (n_3095) );
   NAND2X1 i_550 ( .Y (n_958),
	.B (op_b[31]),
	.A (cmd[1]) );
   OAI21XL i_452 ( .Y (n_955),
	.B0 (n_885),
	.A1 (n_1713),
	.A0 (n_951) );
   NAND2BX1 i_455 ( .Y (n_954),
	.B (op_b[30]),
	.AN (op_a[30]) );
   NOR2BX1 i_542 ( .Y (n_952),
	.B (op_b[30]),
	.AN (op_a[30]) );
   AOI2BB1X1 i_453 ( .Y (n_951),
	.B0 (n_3070),
	.A1N (n_1743),
	.A0N (n_949) );
   AOI21X1 i_454 ( .Y (n_949),
	.B0 (n_1751),
	.A1 (n_1809),
	.A0 (n_1612) );
   OAI211X1 i_436 ( .Y (n_946),
	.C0 (n_945),
	.B0 (n_1762),
	.A1 (n_1766),
	.A0 (n_1765) );
   NAND4BXL i_535 ( .Y (n_945),
	.D (n_1411),
	.C (n_1383),
	.B (n_927),
	.AN (n_1804) );
   OR3XL i_428 ( .Y (n_944),
	.C (n_1213),
	.B (n_1800),
	.A (n_1782) );
   OAI211X1 i_533 ( .Y (n_943),
	.C0 (n_944),
	.B0 (n_1778),
	.A1 (n_1782),
	.A0 (n_1781) );
   NAND2BX1 i_367083 ( .Y (n_942),
	.B (op_b[4]),
	.AN (op_a[4]) );
   NOR2BX1 i_387085 ( .Y (n_940),
	.B (op_a[6]),
	.AN (op_b[6]) );
   NAND2BX1 i_407087 ( .Y (n_937),
	.B (op_b[8]),
	.AN (op_a[8]) );
   NAND2BX1 i_427089 ( .Y (n_935),
	.B (op_b[10]),
	.AN (op_a[10]) );
   NAND2BX1 i_447091 ( .Y (n_933),
	.B (op_b[12]),
	.AN (op_a[12]) );
   NAND2BX1 i_467093 ( .Y (n_931),
	.B (op_b[14]),
	.AN (op_a[14]) );
   NAND2BX1 i_487095 ( .Y (n_929),
	.B (op_b[16]),
	.AN (op_a[16]) );
   NAND2BX1 i_507097 ( .Y (n_927),
	.B (op_b[18]),
	.AN (op_a[18]) );
   NAND2BX1 i_527099 ( .Y (n_925),
	.B (op_b[20]),
	.AN (op_a[20]) );
   NAND2BX1 i_547101 ( .Y (n_923),
	.B (op_b[22]),
	.AN (op_a[22]) );
   NAND2BX1 i_567103 ( .Y (n_921),
	.B (op_b[24]),
	.AN (op_a[24]) );
   OAI21XL i_367 ( .Y (n_917),
	.B0 (n_1812),
	.A1 (n_1703),
	.A0 (n_913) );
   OAI21XL i_514 ( .Y (n_915),
	.B0 (n_917),
	.A1 (op_b[30]),
	.A0 (op_a[30]) );
   AOI21X1 i_368 ( .Y (n_913),
	.B0 (n_1815),
	.A1 (n_3086),
	.A0 (n_1816) );
   AOI211X1 i_369 ( .Y (n_911),
	.C0 (n_909),
	.B0 (n_1819),
	.A1 (n_1823),
	.A0 (n_1822) );
   NOR2X1 i_510 ( .Y (n_909),
	.B (n_1882),
	.A (n_1617) );
   AOI211X1 i_353 ( .Y (n_906),
	.C0 (n_905),
	.B0 (n_1835),
	.A1 (n_1839),
	.A0 (n_1838) );
   NOR4BX1 i_506 ( .Y (n_905),
	.D (n_1416),
	.C (n_1390),
	.B (n_1395),
	.AN (n_1877) );
   NOR4BX1 i_342 ( .Y (n_904),
	.D (n_1218),
	.C (n_1193),
	.B (n_1198),
	.AN (n_1873) );
   AOI211X1 i_504 ( .Y (n_903),
	.C0 (n_904),
	.B0 (n_1851),
	.A1 (n_1855),
	.A0 (n_1854) );
   NAND2BX1 i_937140 ( .Y (n_885),
	.B (op_a[29]),
	.AN (op_b[29]) );
   NAND2BX1 i_412 ( .Y (n_882),
	.B (n_2362),
	.AN (n_2324) );
   NAND2BX1 i_409 ( .Y (n_879),
	.B (n_1758),
	.AN (n_1757) );
   NAND2X1 i_378 ( .Y (n_862),
	.B (n_2062),
	.A (n_2029) );
   NOR2X1 i_377 ( .Y (n_861),
	.B (n_1790),
	.A (n_1789) );
   NAND3X1 i_376 ( .Y (n_860),
	.C (n_3087),
	.B (n_942),
	.A (n_1090) );
   NAND3X1 i_372 ( .Y (n_857),
	.C (n_3065),
	.B (n_1795),
	.A (n_1068) );
   NAND2X1 i_371 ( .Y (n_856),
	.B (n_3065),
	.A (op_a[0]) );
   NOR4BX1 i_332 ( .Y (n_855),
	.D (n_1194),
	.C (n_1100),
	.B (n_1144),
	.AN (n_2103) );
   AOI31X1 i_33 ( .Y (n_828),
	.B0 (n_971),
	.A2 (n_1950),
	.A1 (n_1733),
	.A0 (op_a[31]) );
   NOR2X1 i_9 ( .Y (n_827),
	.B (n_9076575),
	.A (n_1733) );
   AOI22X1 i_1460 ( .Y (n_1620),
	.B1 (n_3069),
	.B0 (n_1640),
	.A1 (n_1716),
	.A0 (n_1613) );
   AOI21X1 i_268 ( .Y (n_1622),
	.B0 (n_1614),
	.A1 (n_1936),
	.A0 (op_a[27]) );
   AOI21X1 i_267 ( .Y (n_1623),
	.B0 (n_1618),
	.A1 (n_911),
	.A0 (n_2382) );
   AND4X1 i_1463 ( .Y (n_1630),
	.D (n_3062),
	.C (n_949),
	.B (n_1640),
	.A (n_3069) );
   NOR4X1 i_1360 ( .Y (n_1632),
	.D (n_1620),
	.C (n_1727),
	.B (n_2387),
	.A (n_1630) );
   OAI21XL i_768552 ( .Y (result[27]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1632) );
   NAND4BXL i_1476 ( .Y (n_1635),
	.D (n_925),
	.C (n_1485),
	.B (n_1534),
	.AN (n_2325) );
   OAI211X1 i_448 ( .Y (n_1637),
	.C0 (n_1635),
	.B0 (n_2324),
	.A1 (n_2325),
	.A0 (n_2294) );
   OAI2BB1X1 i_447 ( .Y (n_1639),
	.B0 (n_2361),
	.A1N (n_2362),
	.A0N (n_1637) );
   NAND2BX1 i_597106 ( .Y (n_1640),
	.B (op_b[27]),
	.AN (op_a[27]) );
   NOR4BX1 i_1485 ( .Y (n_1645),
	.D (n_1541),
	.C (n_1497),
	.B (n_1539),
	.AN (n_2300) );
   NOR2BX1 i_1487 ( .Y (n_1646),
	.B (n_1647),
	.AN (n_2367) );
   AOI211X1 i_363 ( .Y (n_1647),
	.C0 (n_1645),
	.B0 (n_2329),
	.A1 (n_2330),
	.A0 (n_2299) );
   OAI222XL i_1488 ( .Y (n_1648),
	.C1 (n_2366),
	.C0 (n_1646),
	.B1 (op_a[26]),
	.B0 (op_b[26]),
	.A1 (op_a[27]),
	.A0 (op_b[27]) );
   NOR2X1 i_271381 ( .Y (n_1650),
	.B (op_a[27]),
	.A (op_b[27]) );
   NAND2X1 i_1491 ( .Y (n_1652),
	.B (n_2401),
	.A (n_2402) );
   NAND2BX1 i_1496 ( .Y (n_1653),
	.B (n_1654),
	.AN (n_2390) );
   OAI21XL i_275 ( .Y (n_1654),
	.B0 (n_1716),
	.A1 (n_1738),
	.A0 (n_2393) );
   XNOR2X1 i_273 ( .Y (n_1655),
	.B (n_1911),
	.A (op_a[28]) );
   OAI21XL i_272 ( .Y (n_1656),
	.B0 (n_1652),
	.A1 (n_2401),
	.A0 (n_2402) );
   NOR2X1 i_1497 ( .Y (n_1661),
	.B (n_3068),
	.A (n_1655) );
   NAND4BXL i_1369 ( .Y (n_1665),
	.D (n_1653),
	.C (n_2404),
	.B (n_2397),
	.AN (n_1727) );
   OAI2BB1X1 i_758551 ( .Y (result[28]),
	.B0 (n_3060),
	.A1N (n_9076575),
	.A0N (n_1665) );
   AOI31X1 i_449 ( .Y (n_1670),
	.B0 (n_2408),
	.A2 (n_1561),
	.A1 (n_1758),
	.A0 (n_1809) );
   NOR2X1 i_1519 ( .Y (n_1672),
	.B (op_a[29]),
	.A (n_2417) );
   NAND4BXL i_1522 ( .Y (n_1674),
	.D (n_1831),
	.C (n_1881),
	.B (n_1823),
	.AN (n_1567) );
   AOI21X1 i_1525 ( .Y (n_1676),
	.B0 (n_3077),
	.A1 (n_2411),
	.A0 (n_1674) );
   OAI21XL i_1526 ( .Y (n_1678),
	.B0 (n_2413),
	.A1 (n_1815),
	.A0 (n_1676) );
   OAI2BB1X1 i_280 ( .Y (n_1681),
	.B0 (n_1716),
	.A1N (n_3062),
	.A0N (n_2409) );
   AOI21X1 i_279 ( .Y (n_1682),
	.B0 (n_1672),
	.A1 (n_2417),
	.A0 (op_a[29]) );
   OAI31X1 i_278 ( .Y (n_1683),
	.B0 (n_1678),
	.A2 (n_2413),
	.A1 (n_1815),
	.A0 (n_1676) );
   NOR3X1 i_1535 ( .Y (n_1689),
	.C (n_1738),
	.B (n_2406),
	.A (n_2409) );
   AOI211X1 i_1378 ( .Y (n_1692),
	.C0 (n_2423),
	.B0 (n_1727),
	.A1 (n_2406),
	.A0 (n_1681) );
   OAI21XL i_748550 ( .Y (result[29]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1692) );
   NOR4BX1 i_1554 ( .Y (n_1696),
	.D (n_1594),
	.C (n_1497),
	.B (n_1539),
	.AN (n_2367) );
   NOR2X1 i_281382 ( .Y (n_1697),
	.B (op_a[28]),
	.A (op_b[28]) );
   NOR3BX1 i_1557 ( .Y (n_1698),
	.C (n_1699),
	.B (n_1700),
	.AN (n_1816) );
   AOI211X1 i_366 ( .Y (n_1699),
	.C0 (n_1696),
	.B0 (n_2366),
	.A1 (n_2367),
	.A0 (n_2329) );
   NOR2X1 i_261380 ( .Y (n_1700),
	.B (op_a[26]),
	.A (op_b[26]) );
   NOR2X1 i_291383 ( .Y (n_1703),
	.B (op_a[29]),
	.A (op_b[29]) );
   AOI221X1 i_365 ( .Y (n_1704),
	.C0 (n_1698),
	.B1 (op_b[28]),
	.B0 (op_a[28]),
	.A1 (n_3066),
	.A0 (n_2399) );
   NAND3BX1 i_1561 ( .Y (n_1705),
	.C (n_1587),
	.B (n_2362),
	.AN (n_2325) );
   NAND2BX1 i_607107 ( .Y (n_1706),
	.B (op_b[28]),
	.AN (op_a[28]) );
   NAND3X1 i_451 ( .Y (n_1708),
	.C (n_1705),
	.B (n_2361),
	.A (n_882) );
   NAND2BX1 i_587105 ( .Y (n_1709),
	.B (op_b[26]),
	.AN (op_a[26]) );
   NOR2BX1 i_927139 ( .Y (n_1710),
	.B (op_b[28]),
	.AN (op_a[28]) );
   NOR2BX1 i_617108 ( .Y (n_1713),
	.B (op_a[29]),
	.AN (op_b[29]) );
   AOI221X1 i_450 ( .Y (n_1714),
	.C0 (n_1710),
	.B1 (n_2426),
	.B0 (n_1708),
	.A1 (n_1706),
	.A0 (n_2391) );
   NAND3BX1 i_1092 ( .Y (n_1716),
	.C (n_1736),
	.B (cmd[2]),
	.AN (cmd[0]) );
   OAI21XL i_288 ( .Y (n_1720),
	.B0 (n_2436),
	.A1 (n_3068),
	.A0 (n_2434) );
   OAI221XL i_2879002 ( .Y (n_1722),
	.C0 (n_1716),
	.B1 (n_3088),
	.B0 (n_1738),
	.A1 (n_3095),
	.A0 (n_2431) );
   AOI22X1 i_285 ( .Y (n_1723),
	.B1 (n_868),
	.B0 (n_2431),
	.A1 (n_3062),
	.A0 (n_3088) );
   NOR2X1 i_10 ( .Y (n_1727),
	.B (n_3068),
	.A (n_1915) );
   AOI21X1 i_1387 ( .Y (n_1730),
	.B0 (n_2441),
	.A1 (n_2425),
	.A0 (n_1722) );
   OAI21XL i_738549 ( .Y (result[30]),
	.B0 (n_3060),
	.A1 (n_907),
	.A0 (n_1730) );
   AOI21X1 i_1396 ( .Y (n_1733),
	.B0 (n_1949),
	.A1 (n_1740),
	.A0 (n_962) );
   NAND2X1 i_1587 ( .Y (n_1734),
	.B (n_907),
	.A (n_1733) );
   OAI21XL i_728548 ( .Y (result[31]),
	.B0 (n_1734),
	.A1 (n_907),
	.A0 (n_1733) );
   NOR2X1 i_14 ( .Y (n_1736),
	.B (cmd[1]),
	.A (cmd[3]) );
   NAND3BX1 i_1081 ( .Y (n_1738),
	.C (n_1736),
	.B (cmd[0]),
	.AN (cmd[2]) );
   XOR2X1 i_1607206 ( .Y (n_1740),
	.B (op_b[31]),
	.A (op_a[31]) );
   NOR2BX1 i_917138 ( .Y (n_1741),
	.B (op_b[27]),
	.AN (op_a[27]) );
   AOI21X1 i_1897235 ( .Y (n_1742),
	.B0 (n_1710),
	.A1 (n_1741),
	.A0 (n_1706) );
   NAND2X1 i_13 ( .Y (n_1743),
	.B (n_1640),
	.A (n_1706) );
   NOR2BX1 i_907137 ( .Y (n_1744),
	.B (op_b[26]),
	.AN (op_a[26]) );
   NOR2BX1 i_897136 ( .Y (n_1745),
	.B (op_b[25]),
	.AN (op_a[25]) );
   AOI21X1 i_1877233 ( .Y (n_1746),
	.B0 (n_1744),
	.A1 (n_1745),
	.A0 (n_1709) );
   NOR2BX1 i_887135 ( .Y (n_1747),
	.B (op_b[24]),
	.AN (op_a[24]) );
   NOR2BX1 i_877134 ( .Y (n_1748),
	.B (op_b[23]),
	.AN (op_a[23]) );
   AOI21X1 i_1857231 ( .Y (n_1749),
	.B0 (n_1747),
	.A1 (n_1748),
	.A0 (n_921) );
   NAND2X1 i_2197263 ( .Y (n_1750),
	.B (n_1585),
	.A (n_1709) );
   OAI21XL i_2507290 ( .Y (n_1751),
	.B0 (n_1746),
	.A1 (n_1749),
	.A0 (n_1750) );
   NOR2BX1 i_867133 ( .Y (n_1752),
	.B (op_b[22]),
	.AN (op_a[22]) );
   NOR2BX1 i_857132 ( .Y (n_1753),
	.B (op_b[21]),
	.AN (op_a[21]) );
   AOI21X1 i_1837229 ( .Y (n_1754),
	.B0 (n_1752),
	.A1 (n_1753),
	.A0 (n_923) );
   NOR2BX1 i_847131 ( .Y (n_1755),
	.B (op_b[20]),
	.AN (op_a[20]) );
   NOR2BX1 i_837130 ( .Y (n_1756),
	.B (op_b[19]),
	.AN (op_a[19]) );
   AOI21X1 i_1817227 ( .Y (n_1757),
	.B0 (n_1755),
	.A1 (n_1756),
	.A0 (n_925) );
   AND2X1 i_2157259 ( .Y (n_1758),
	.B (n_1485),
	.A (n_923) );
   NOR2BX1 i_827129 ( .Y (n_1760),
	.B (op_b[18]),
	.AN (op_a[18]) );
   NOR2BX1 i_817128 ( .Y (n_1761),
	.B (op_b[17]),
	.AN (op_a[17]) );
   AOI21X1 i_1797225 ( .Y (n_1762),
	.B0 (n_1760),
	.A1 (n_1761),
	.A0 (n_927) );
   NOR2BX1 i_807127 ( .Y (n_1763),
	.B (op_b[16]),
	.AN (op_a[16]) );
   NOR2BX1 i_797126 ( .Y (n_1764),
	.B (op_b[15]),
	.AN (op_a[15]) );
   AOI21X1 i_1777223 ( .Y (n_1765),
	.B0 (n_1763),
	.A1 (n_1764),
	.A0 (n_929) );
   NAND2X1 i_2117255 ( .Y (n_1766),
	.B (n_1383),
	.A (n_927) );
   NOR2BX1 i_787125 ( .Y (n_1768),
	.B (op_b[14]),
	.AN (op_a[14]) );
   NOR2BX1 i_777124 ( .Y (n_1769),
	.B (op_b[13]),
	.AN (op_a[13]) );
   AOI21X1 i_1757221 ( .Y (n_1770),
	.B0 (n_1768),
	.A1 (n_1769),
	.A0 (n_931) );
   NOR2BX1 i_767123 ( .Y (n_1771),
	.B (op_b[12]),
	.AN (op_a[12]) );
   NOR2BX1 i_757122 ( .Y (n_1772),
	.B (op_b[11]),
	.AN (op_a[11]) );
   AOI21X1 i_1737219 ( .Y (n_1773),
	.B0 (n_1771),
	.A1 (n_1772),
	.A0 (n_933) );
   NAND2X1 i_2077251 ( .Y (n_1774),
	.B (n_1286),
	.A (n_931) );
   NOR2BX1 i_747121 ( .Y (n_1776),
	.B (op_b[10]),
	.AN (op_a[10]) );
   NOR2BX1 i_737120 ( .Y (n_1777),
	.B (op_b[9]),
	.AN (op_a[9]) );
   AOI21X1 i_1717217 ( .Y (n_1778),
	.B0 (n_1776),
	.A1 (n_1777),
	.A0 (n_935) );
   NOR2BX1 i_727119 ( .Y (n_1779),
	.B (op_b[8]),
	.AN (op_a[8]) );
   NOR2BX1 i_717118 ( .Y (n_1780),
	.B (op_b[7]),
	.AN (op_a[7]) );
   AOI21X1 i_1697215 ( .Y (n_1781),
	.B0 (n_1779),
	.A1 (n_1780),
	.A0 (n_937) );
   NAND2X1 i_2037247 ( .Y (n_1782),
	.B (n_1186),
	.A (n_935) );
   NOR2BX1 i_707117 ( .Y (n_1784),
	.B (op_b[6]),
	.AN (op_a[6]) );
   NAND2BX1 i_697116 ( .Y (n_1785),
	.B (op_a[5]),
	.AN (op_b[5]) );
   OAI21XL i_1677213 ( .Y (n_1786),
	.B0 (n_3074),
	.A1 (n_940),
	.A0 (n_1785) );
   NOR2BX1 i_687115 ( .Y (n_1787),
	.B (op_b[4]),
	.AN (op_a[4]) );
   NOR2BX1 i_677114 ( .Y (n_1788),
	.B (op_b[3]),
	.AN (op_a[3]) );
   AOI21X1 i_1657211 ( .Y (n_1789),
	.B0 (n_1787),
	.A1 (n_1788),
	.A0 (n_942) );
   NAND2BX1 i_1997243 ( .Y (n_1790),
	.B (n_1090),
	.AN (n_940) );
   NOR2BX1 i_667113 ( .Y (n_1792),
	.B (op_b[2]),
	.AN (op_a[2]) );
   NOR2BX1 i_657112 ( .Y (n_1793),
	.B (op_b[1]),
	.AN (op_a[1]) );
   AOI21X1 i_1637209 ( .Y (n_1794),
	.B0 (n_1792),
	.A1 (n_1793),
	.A0 (n_1068) );
   NAND2BX1 i_1617207 ( .Y (n_1795),
	.B (op_b[0]),
	.AN (op_a[0]) );
   NAND2X1 i_2267266 ( .Y (n_1797),
	.B (n_1794),
	.A (n_857) );
   NAND2X1 i_1977241 ( .Y (n_1798),
	.B (n_1045),
	.A (n_942) );
   NOR2X1 i_531 ( .Y (n_1799),
	.B (n_1798),
	.A (n_1790) );
   NAND2X1 i_2017245 ( .Y (n_1800),
	.B (n_1135),
	.A (n_937) );
   NAND2X1 i_2057249 ( .Y (n_1802),
	.B (n_1237),
	.A (n_933) );
   NAND2X1 i_2097253 ( .Y (n_1804),
	.B (n_1332),
	.A (n_929) );
   NAND2X1 i_2137257 ( .Y (n_1806),
	.B (n_1434),
	.A (n_925) );
   NAND2X1 i_2177261 ( .Y (n_1808),
	.B (n_1532),
	.A (n_921) );
   NOR2X1 i_15 ( .Y (n_1809),
	.B (n_1808),
	.A (n_1750) );
   AOI21X1 i_443 ( .Y (n_1810),
	.B0 (n_952),
	.A1 (n_954),
	.A0 (n_955) );
   NAND2X1 i_611415 ( .Y (n_1812),
	.B (op_b[29]),
	.A (op_a[29]) );
   NAND2X1 i_601414 ( .Y (n_1813),
	.B (op_b[28]),
	.A (op_a[28]) );
   NAND2X1 i_591413 ( .Y (n_1814),
	.B (op_b[27]),
	.A (op_a[27]) );
   OAI21XL i_1561510 ( .Y (n_1815),
	.B0 (n_1813),
	.A1 (n_1697),
	.A0 (n_1814) );
   NOR2X1 i_12 ( .Y (n_1816),
	.B (n_1697),
	.A (n_1650) );
   NAND2X1 i_581412 ( .Y (n_1817),
	.B (op_b[26]),
	.A (op_a[26]) );
   NAND2X1 i_571411 ( .Y (n_1818),
	.B (op_b[25]),
	.A (op_a[25]) );
   OAI21XL i_1541508 ( .Y (n_1819),
	.B0 (n_1817),
	.A1 (n_1818),
	.A0 (n_1700) );
   NAND2X1 i_561410 ( .Y (n_1820),
	.B (op_b[24]),
	.A (op_a[24]) );
   NAND2X1 i_551409 ( .Y (n_1821),
	.B (op_b[23]),
	.A (op_a[23]) );
   OAI21XL i_1521506 ( .Y (n_1822),
	.B0 (n_1820),
	.A1 (n_1821),
	.A0 (n_1544) );
   NOR2X1 i_185 ( .Y (n_1823),
	.B (n_1592),
	.A (n_1700) );
   NAND2X1 i_541408 ( .Y (n_1825),
	.B (op_b[22]),
	.A (op_a[22]) );
   NAND2X1 i_531407 ( .Y (n_1826),
	.B (op_b[21]),
	.A (op_a[21]) );
   OAI21XL i_1501504 ( .Y (n_1827),
	.B0 (n_1825),
	.A1 (n_1826),
	.A0 (n_1497) );
   NAND2X1 i_521406 ( .Y (n_1828),
	.B (op_b[20]),
	.A (op_a[20]) );
   NAND2X1 i_511405 ( .Y (n_1829),
	.B (op_b[19]),
	.A (op_a[19]) );
   OAI21XL i_1481502 ( .Y (n_1830),
	.B0 (n_1828),
	.A1 (n_1829),
	.A0 (n_1446) );
   NOR2X1 i_181 ( .Y (n_1831),
	.B (n_1492),
	.A (n_1497) );
   NAND2X1 i_501404 ( .Y (n_1833),
	.B (op_b[18]),
	.A (op_a[18]) );
   NAND2X1 i_491403 ( .Y (n_1834),
	.B (op_b[17]),
	.A (op_a[17]) );
   OAI21XL i_1461500 ( .Y (n_1835),
	.B0 (n_1833),
	.A1 (n_1834),
	.A0 (n_1395) );
   NAND2X1 i_481402 ( .Y (n_1836),
	.B (op_b[16]),
	.A (op_a[16]) );
   NAND2X1 i_471401 ( .Y (n_1837),
	.B (op_b[15]),
	.A (op_a[15]) );
   OAI21XL i_1441498 ( .Y (n_1838),
	.B0 (n_1836),
	.A1 (n_1837),
	.A0 (n_1344) );
   NOR2X1 i_177 ( .Y (n_1839),
	.B (n_1390),
	.A (n_1395) );
   NAND2X1 i_461400 ( .Y (n_1841),
	.B (op_b[14]),
	.A (op_a[14]) );
   NAND2X1 i_451399 ( .Y (n_1842),
	.B (op_b[13]),
	.A (op_a[13]) );
   OAI21XL i_1421496 ( .Y (n_1843),
	.B0 (n_1841),
	.A1 (n_1842),
	.A0 (n_1297) );
   NAND2X1 i_441398 ( .Y (n_1844),
	.B (op_b[12]),
	.A (op_a[12]) );
   NAND2X1 i_431397 ( .Y (n_1845),
	.B (op_b[11]),
	.A (op_a[11]) );
   OAI21XL i_1401494 ( .Y (n_1846),
	.B0 (n_1844),
	.A1 (n_1845),
	.A0 (n_1249) );
   NOR2X1 i_173 ( .Y (n_1847),
	.B (n_1293),
	.A (n_1297) );
   NAND2X1 i_421396 ( .Y (n_1849),
	.B (op_b[10]),
	.A (op_a[10]) );
   NAND2X1 i_411395 ( .Y (n_1850),
	.B (op_b[9]),
	.A (op_a[9]) );
   OAI21XL i_1381492 ( .Y (n_1851),
	.B0 (n_1849),
	.A1 (n_1850),
	.A0 (n_1198) );
   NAND2X1 i_401394 ( .Y (n_1852),
	.B (op_b[8]),
	.A (op_a[8]) );
   NAND2X1 i_391393 ( .Y (n_1853),
	.B (op_b[7]),
	.A (op_a[7]) );
   OAI21XL i_1361490 ( .Y (n_1854),
	.B0 (n_1852),
	.A1 (n_1853),
	.A0 (n_1147) );
   NOR2X1 i_169 ( .Y (n_1855),
	.B (n_1193),
	.A (n_1198) );
   NAND2X1 i_381392 ( .Y (n_1857),
	.B (op_b[6]),
	.A (op_a[6]) );
   NAND2X1 i_371391 ( .Y (n_1858),
	.B (op_b[5]),
	.A (op_a[5]) );
   OAI21XL i_1341488 ( .Y (n_1859),
	.B0 (n_1857),
	.A1 (n_1858),
	.A0 (n_1100) );
   NAND2X1 i_361390 ( .Y (n_1860),
	.B (op_b[4]),
	.A (op_a[4]) );
   NAND2X1 i_351389 ( .Y (n_1861),
	.B (op_b[3]),
	.A (op_a[3]) );
   OAI21XL i_1321486 ( .Y (n_1862),
	.B0 (n_1860),
	.A1 (n_1861),
	.A0 (n_1053) );
   NOR2X1 i_1651517 ( .Y (n_1863),
	.B (n_1095),
	.A (n_1100) );
   NAND2X1 i_341388 ( .Y (n_1865),
	.B (op_b[2]),
	.A (op_a[2]) );
   NAND2X1 i_331387 ( .Y (n_1866),
	.B (op_b[1]),
	.A (op_a[1]) );
   OAI21XL i_1301484 ( .Y (n_1867),
	.B0 (n_1865),
	.A1 (n_1866),
	.A0 (n_1096) );
   NAND2X1 i_321386 ( .Y (n_1868),
	.B (op_b[0]),
	.A (op_a[0]) );
   NOR2X1 i_498 ( .Y (n_1869),
	.B (n_1072),
	.A (n_1096) );
   AOI21X1 i_192 ( .Y (n_1870),
	.B0 (n_1867),
	.A1 (n_3085),
	.A0 (n_1869) );
   NOR2X1 i_1631515 ( .Y (n_1871),
	.B (n_1097),
	.A (n_1053) );
   NOR2X1 i_1671519 ( .Y (n_1873),
	.B (n_1144),
	.A (n_1147) );
   NOR2X1 i_171 ( .Y (n_1875),
	.B (n_1244),
	.A (n_1249) );
   NOR2X1 i_175 ( .Y (n_1877),
	.B (n_1339),
	.A (n_1344) );
   NOR2X1 i_179 ( .Y (n_1879),
	.B (n_1441),
	.A (n_1446) );
   NAND2X1 i_509 ( .Y (n_1880),
	.B (n_1879),
	.A (n_1831) );
   NOR2X1 i_183 ( .Y (n_1881),
	.B (n_1539),
	.A (n_1544) );
   NAND2X1 i_16 ( .Y (n_1882),
	.B (n_1881),
	.A (n_1823) );
   OAI2BB1X1 i_406 ( .Y (n_1883),
	.B0 (n_915),
	.A1N (op_b[30]),
	.A0N (op_a[30]) );
   NOR2X1 i_11787 ( .Y (n_1885),
	.B (op_a[1]),
	.A (op_a[0]) );
   NOR3X1 i_341819 ( .Y (n_1886),
	.C (op_a[2]),
	.B (op_a[1]),
	.A (op_a[0]) );
   NOR2X1 i_26 ( .Y (n_1887),
	.B (op_a[7]),
	.A (op_a[6]) );
   NOR2X1 i_25 ( .Y (n_1888),
	.B (op_a[5]),
	.A (op_a[4]) );
   NAND4BXL i_711854 ( .Y (n_1891),
	.D (n_1886),
	.C (n_1887),
	.B (n_1888),
	.AN (op_a[3]) );
   NOR2X1 i_27 ( .Y (n_1892),
	.B (op_a[9]),
	.A (op_a[8]) );
   NOR2X1 i_28 ( .Y (n_1893),
	.B (op_a[11]),
	.A (op_a[10]) );
   NAND3BX1 i_1071887 ( .Y (n_1895),
	.C (n_1893),
	.B (n_1892),
	.AN (n_1891) );
   NOR2X1 i_30 ( .Y (n_1896),
	.B (op_a[14]),
	.A (op_a[13]) );
   NOR4BX1 i_1111891 ( .Y (n_1899),
	.D (n_1895),
	.C (op_a[15]),
	.B (op_a[12]),
	.AN (n_1896) );
   NOR2X1 i_24 ( .Y (n_1900),
	.B (op_a[17]),
	.A (op_a[16]) );
   NOR2X1 i_31 ( .Y (n_1901),
	.B (op_a[19]),
	.A (op_a[18]) );
   NAND3X1 i_1471921 ( .Y (n_1903),
	.C (n_1899),
	.B (n_1901),
	.A (n_1900) );
   NOR2X1 i_29 ( .Y (n_1904),
	.B (op_a[23]),
	.A (op_a[22]) );
   NOR2X1 i_32 ( .Y (n_1905),
	.B (op_a[21]),
	.A (op_a[20]) );
   NOR4BX1 i_1511925 ( .Y (n_1907),
	.D (n_1903),
	.C (op_a[21]),
	.B (op_a[20]),
	.AN (n_1904) );
   NOR2X1 i_20 ( .Y (n_1908),
	.B (op_a[27]),
	.A (op_a[26]) );
   NOR2X1 i_21 ( .Y (n_1909),
	.B (op_a[25]),
	.A (op_a[24]) );
   NAND3X1 i_1551929 ( .Y (n_1911),
	.C (n_1907),
	.B (n_1908),
	.A (n_1909) );
   NOR2X1 i_22 ( .Y (n_1912),
	.B (op_a[29]),
	.A (op_a[28]) );
   NAND2X1 i_8 ( .Y (n_1915),
	.B (n_166),
	.A (ovm) );
   NAND3X1 i_1095 ( .Y (n_1917),
	.C (n_1736),
	.B (cmd[2]),
	.A (cmd[0]) );
   NOR2BX1 i_3 ( .Y (n_1918),
	.B (n_1917),
	.AN (op_a[31]) );
   NOR2X1 i_459 ( .Y (n_1919),
	.B (op_a[6]),
	.A (op_a[3]) );
   NAND3X1 i_701853 ( .Y (n_1921),
	.C (n_1886),
	.B (n_1888),
	.A (n_1919) );
   NOR4BX1 i_1061886 ( .Y (n_1924),
	.D (n_1921),
	.C (op_a[10]),
	.B (op_a[7]),
	.AN (n_1892) );
   NOR4X1 i_464 ( .Y (n_1926),
	.D (op_a[14]),
	.C (op_a[13]),
	.B (op_a[12]),
	.A (op_a[11]) );
   NAND2X1 i_1101890 ( .Y (n_1927),
	.B (n_1924),
	.A (n_1926) );
   NOR4BX1 i_1461920 ( .Y (n_1930),
	.D (n_1927),
	.C (op_a[18]),
	.B (op_a[15]),
	.AN (n_1900) );
   NOR4X1 i_468 ( .Y (n_1932),
	.D (op_a[21]),
	.C (op_a[20]),
	.B (op_a[22]),
	.A (op_a[19]) );
   NAND2X1 i_1501924 ( .Y (n_1933),
	.B (n_1930),
	.A (n_1932) );
   NOR4BX1 i_1541928 ( .Y (n_1936),
	.D (n_1933),
	.C (op_a[26]),
	.B (op_a[23]),
	.AN (n_1909) );
   NOR4X1 i_561 ( .Y (n_1938),
	.D (op_a[29]),
	.C (op_a[28]),
	.B (op_a[30]),
	.A (op_a[27]) );
   NAND3BX1 i_1088 ( .Y (n_1942),
	.C (cmd[0]),
	.B (cmd[1]),
	.AN (cmd[2]) );
   NAND3BX1 i_1098 ( .Y (n_1944),
	.C (cmd[1]),
	.B (cmd[2]),
	.AN (cmd[0]) );
   AND2X1 i_1100 ( .Y (n_1946),
	.B (cmd[1]),
	.A (cmd[0]) );
   AOI22X1 i_564 ( .Y (n_1947),
	.B1 (op_a[31]),
	.B0 (n_963),
	.A1 (n_1946),
	.A0 (op_b[31]) );
   OAI211X1 i_566 ( .Y (n_1949),
	.C0 (n_1947),
	.B0 (n_967),
	.A1 (n_1740),
	.A0 (n_964) );
   AOI21X1 i_11 ( .Y (n_1950),
	.B0 (n_970),
	.A1 (n_3095),
	.A0 (op_b[31]) );
   NAND4BXL i_578 ( .Y (n_1955),
	.D (n_1942),
	.C (n_1917),
	.B (n_1944),
	.AN (n_974) );
   AOI221X1 i_586 ( .Y (n_1957),
	.C0 (n_1727),
	.B1 (n_3085),
	.B0 (cmd[1]),
	.A1 (op_b[0]),
	.A0 (n_978) );
   NAND2X1 i_39 ( .Y (n_1959),
	.B (n_3065),
	.A (n_3075) );
   NAND2X1 i_42 ( .Y (n_1961),
	.B (op_a[0]),
	.A (op_a[31]) );
   AOI21X1 i_593 ( .Y (n_1962),
	.B0 (n_986),
	.A1 (op_a[1]),
	.A0 (n_1961) );
   AOI222X1 i_607 ( .Y (n_1965),
	.C1 (op_b[1]),
	.C0 (n_1946),
	.B1 (n_3063),
	.B0 (op_a[1]),
	.A1 (n_3083),
	.A0 (cmd[1]) );
   OAI21XL i_608 ( .Y (n_1966),
	.B0 (n_1965),
	.A1 (n_1942),
	.A0 (n_1072) );
   AOI211X1 i_610 ( .Y (n_1968),
	.C0 (n_999),
	.B0 (n_1966),
	.A1 (n_868),
	.A0 (n_993) );
   OAI31X1 i_611 ( .Y (n_1969),
	.B0 (n_1968),
	.A2 (n_1738),
	.A1 (n_1795),
	.A0 (n_1959) );
   NAND2BX1 i_45 ( .Y (n_1970),
	.B (n_1068),
	.AN (n_1792) );
   OAI21XL i_1627208 ( .Y (n_1971),
	.B0 (n_3075),
	.A1 (n_1136),
	.A0 (op_b[0]) );
   NAND2BX1 i_2257265 ( .Y (n_1972),
	.B (n_856),
	.AN (n_1971) );
   OAI21XL i_48 ( .Y (n_1974),
	.B0 (op_a[31]),
	.A1 (op_a[1]),
	.A0 (op_a[0]) );
   AOI21X1 i_618 ( .Y (n_1975),
	.B0 (n_1006),
	.A1 (op_a[2]),
	.A0 (n_1974) );
   OAI21XL i_1291483 ( .Y (n_1976),
	.B0 (n_1866),
	.A1 (n_1868),
	.A0 (n_1072) );
   NOR2X1 i_47 ( .Y (n_1977),
	.B (n_3084),
	.A (n_1096) );
   AOI222X1 i_633 ( .Y (n_1979),
	.C1 (op_b[2]),
	.C0 (n_1946),
	.B1 (n_3063),
	.B0 (op_a[2]),
	.A1 (n_3084),
	.A0 (cmd[1]) );
   OAI21XL i_634 ( .Y (n_1980),
	.B0 (n_1979),
	.A1 (n_1942),
	.A0 (n_1096) );
   AOI211X1 i_636 ( .Y (n_1982),
	.C0 (n_1020),
	.B0 (n_1980),
	.A1 (n_868),
	.A0 (n_1014) );
   OAI31X1 i_637 ( .Y (n_1983),
	.B0 (n_1982),
	.A2 (n_1972),
	.A1 (n_1738),
	.A0 (n_1970) );
   NAND2BX1 i_51 ( .Y (n_1984),
	.B (n_1045),
	.AN (n_1788) );
   NAND2X1 i_54 ( .Y (n_1986),
	.B (n_3067),
	.A (op_a[31]) );
   AOI21X1 i_643 ( .Y (n_1987),
	.B0 (n_1026),
	.A1 (n_1986),
	.A0 (op_a[3]) );
   NOR2X1 i_53 ( .Y (n_1988),
	.B (n_3081),
	.A (n_1097) );
   AOI222X1 i_657 ( .Y (n_1990),
	.C1 (op_b[3]),
	.C0 (n_1946),
	.B1 (n_3063),
	.B0 (op_a[3]),
	.A1 (n_3081),
	.A0 (cmd[1]) );
   OAI21XL i_658 ( .Y (n_1991),
	.B0 (n_1990),
	.A1 (n_1942),
	.A0 (n_1097) );
   AOI211X1 i_660 ( .Y (n_1993),
	.C0 (n_1039),
	.B0 (n_1991),
	.A1 (n_868),
	.A0 (n_1033) );
   OAI31X1 i_661 ( .Y (n_1994),
	.B0 (n_1993),
	.A2 (n_1738),
	.A1 (n_1797),
	.A0 (n_1984) );
   NAND2BX1 i_57 ( .Y (n_1995),
	.B (n_942),
	.AN (n_1787) );
   AOI21X1 i_1647210 ( .Y (n_1996),
	.B0 (n_1788),
	.A1 (n_1792),
	.A0 (n_1045) );
   NAND2X1 i_1967240 ( .Y (n_1997),
	.B (n_1068),
	.A (n_1045) );
   AOI31X1 i_2277267 ( .Y (n_1998),
	.B0 (n_3087),
	.A2 (n_1068),
	.A1 (n_1045),
	.A0 (n_1971) );
   OAI21XL i_17 ( .Y (n_2000),
	.B0 (op_a[31]),
	.A1 (n_3067),
	.A0 (op_a[3]) );
   AOI21X1 i_671 ( .Y (n_2001),
	.B0 (n_1048),
	.A1 (op_a[4]),
	.A0 (n_2000) );
   OAI21XL i_1311485 ( .Y (n_2002),
	.B0 (n_1861),
	.A1 (n_1865),
	.A0 (n_1097) );
   NOR2X1 i_674 ( .Y (n_2003),
	.B (n_1096),
	.A (n_1097) );
   AOI21X1 i_193 ( .Y (n_2004),
	.B0 (n_2002),
	.A1 (n_2003),
	.A0 (n_1976) );
   NOR2X1 i_59 ( .Y (n_2005),
	.B (n_3082),
	.A (n_1053) );
   AOI222X1 i_687 ( .Y (n_2007),
	.C1 (op_b[4]),
	.C0 (n_1946),
	.B1 (n_3063),
	.B0 (op_a[4]),
	.A1 (n_3082),
	.A0 (cmd[1]) );
   OAI21XL i_688 ( .Y (n_2008),
	.B0 (n_2007),
	.A1 (n_1942),
	.A0 (n_1053) );
   AOI211X1 i_690 ( .Y (n_2010),
	.C0 (n_1063),
	.B0 (n_2008),
	.A1 (n_868),
	.A0 (n_1057) );
   OAI31X1 i_691 ( .Y (n_2011),
	.B0 (n_2010),
	.A2 (n_1738),
	.A1 (n_1995),
	.A0 (n_1137) );
   OAI21XL i_2287268 ( .Y (n_2013),
	.B0 (n_1789),
	.A1 (n_1794),
	.A0 (n_1798) );
   NOR2X1 i_699 ( .Y (n_2016),
	.B (op_a[3]),
	.A (op_a[2]) );
   NOR4BX1 i_681851 ( .Y (n_2017),
	.D (op_a[4]),
	.C (op_a[3]),
	.B (op_a[2]),
	.AN (n_1885) );
   NAND2BX1 i_65 ( .Y (n_2018),
	.B (op_a[31]),
	.AN (n_2017) );
   AOI21X1 i_702 ( .Y (n_2019),
	.B0 (n_1070),
	.A1 (n_2018),
	.A0 (op_a[5]) );
   AOI21X1 i_194 ( .Y (n_2020),
	.B0 (n_1862),
	.A1 (n_1871),
	.A0 (n_1867) );
   NOR2X1 i_64 ( .Y (n_2021),
	.B (n_3079),
	.A (n_1095) );
   AOI222X1 i_718 ( .Y (n_2023),
	.C1 (op_b[5]),
	.C0 (n_1946),
	.B1 (n_3063),
	.B0 (op_a[5]),
	.A1 (n_3079),
	.A0 (cmd[1]) );
   OAI221XL i_720 ( .Y (n_2025),
	.C0 (n_2023),
	.B1 (n_3095),
	.B0 (n_1078),
	.A1 (n_1942),
	.A0 (n_1095) );
   NAND2BX1 i_68 ( .Y (n_2028),
	.B (n_3074),
	.AN (n_940) );
   NAND2X1 i_1667212 ( .Y (n_2029),
	.B (n_1785),
	.A (n_1089) );
   NAND3X1 i_691852 ( .Y (n_2035),
	.C (n_1885),
	.B (n_2016),
	.A (n_1888) );
   NAND2X1 i_72 ( .Y (n_2036),
	.B (op_a[31]),
	.A (n_2035) );
   AOI21X1 i_733 ( .Y (n_2037),
	.B0 (n_1092),
	.A1 (op_a[6]),
	.A0 (n_2036) );
   OAI21XL i_1331487 ( .Y (n_2038),
	.B0 (n_1858),
	.A1 (n_1860),
	.A0 (n_1095) );
   NOR2X1 i_1641516 ( .Y (n_2039),
	.B (n_1053),
	.A (n_1095) );
   AOI21X1 i_195 ( .Y (n_2040),
	.B0 (n_2038),
	.A1 (n_2039),
	.A0 (n_2002) );
   NOR2X1 i_70 ( .Y (n_2042),
	.B (n_3080),
	.A (n_1100) );
   AOI222X1 i_750 ( .Y (n_2044),
	.C1 (op_b[6]),
	.C0 (n_1946),
	.B1 (n_3063),
	.B0 (op_a[6]),
	.A1 (n_3080),
	.A0 (cmd[1]) );
   OAI21XL i_751 ( .Y (n_2045),
	.B0 (n_2044),
	.A1 (n_1942),
	.A0 (n_1100) );
   AOI211X1 i_753 ( .Y (n_2047),
	.C0 (n_1110),
	.B0 (n_2045),
	.A1 (n_868),
	.A0 (n_1104) );
   OAI31X1 i_754 ( .Y (n_2048),
	.B0 (n_2047),
	.A2 (n_1187),
	.A1 (n_1738),
	.A0 (n_2028) );
   NAND2BX1 i_75 ( .Y (n_2049),
	.B (n_1135),
	.AN (n_1780) );
   NAND2X1 i_78 ( .Y (n_2051),
	.B (op_a[31]),
	.A (n_1921) );
   AOI21X1 i_760 ( .Y (n_2052),
	.B0 (n_1116),
	.A1 (op_a[7]),
	.A0 (n_2051) );
   NOR2X1 i_77 ( .Y (n_2053),
	.B (n_3078),
	.A (n_1144) );
   AOI222X1 i_774 ( .Y (n_2055),
	.C1 (op_b[7]),
	.C0 (n_1946),
	.B1 (n_3063),
	.B0 (op_a[7]),
	.A1 (n_3078),
	.A0 (cmd[1]) );
   OAI21XL i_775 ( .Y (n_2056),
	.B0 (n_2055),
	.A1 (n_1942),
	.A0 (n_1144) );
   AOI211X1 i_777 ( .Y (n_2058),
	.C0 (n_1129),
	.B0 (n_2056),
	.A1 (n_868),
	.A0 (n_1123) );
   OAI31X1 i_778 ( .Y (n_2059),
	.B0 (n_2058),
	.A2 (n_3076),
	.A1 (n_1738),
	.A0 (n_2049) );
   NAND2BX1 i_82 ( .Y (n_2060),
	.B (n_937),
	.AN (n_1779) );
   AOI21X1 i_1687214 ( .Y (n_2061),
	.B0 (n_1780),
	.A1 (n_1784),
	.A0 (n_1135) );
   NOR2BX1 i_2007244 ( .Y (n_2062),
	.B (n_940),
	.AN (n_1135) );
   OAI21XL i_1351489 ( .Y (n_2066),
	.B0 (n_1853),
	.A1 (n_1857),
	.A0 (n_1144) );
   NOR2X1 i_1661518 ( .Y (n_2067),
	.B (n_1100),
	.A (n_1144) );
   AOI21X1 i_83 ( .Y (n_2070),
	.B0 (n_1147),
	.A1 (op_b[8]),
	.A0 (op_a[8]) );
   OAI21XL i_0 ( .Y (n_2071),
	.B0 (n_1944),
	.A1 (n_1917),
	.A0 (op_a[31]) );
   OAI211X1 i_804 ( .Y (n_2072),
	.C0 (cmd[1]),
	.B0 (op_b[8]),
	.A1 (cmd[0]),
	.A0 (op_a[8]) );
   OAI221XL i_806 ( .Y (n_2074),
	.C0 (n_2072),
	.B1 (n_3068),
	.B0 (n_1150),
	.A1 (n_1942),
	.A0 (n_1147) );
   AOI221X1 i_808 ( .Y (n_2076),
	.C0 (n_2074),
	.B1 (n_868),
	.B0 (n_1151),
	.A1 (op_a[8]),
	.A0 (n_2071) );
   OAI31X1 i_809 ( .Y (n_2077),
	.B0 (n_2076),
	.A2 (n_1238),
	.A1 (n_1738),
	.A0 (n_2060) );
   NAND2BX1 i_87 ( .Y (n_2079),
	.B (n_1186),
	.AN (n_1777) );
   AOI31X1 i_2327272 ( .Y (n_2080),
	.B0 (n_3073),
	.A2 (n_1135),
	.A1 (n_1786),
	.A0 (n_937) );
   AOI21X1 i_198 ( .Y (n_2083),
	.B0 (n_1854),
	.A1 (n_1873),
	.A0 (n_1859) );
   AOI21X1 i_88 ( .Y (n_2085),
	.B0 (n_1193),
	.A1 (op_b[9]),
	.A0 (op_a[9]) );
   NOR4X1 i_818 ( .Y (n_2087),
	.D (op_a[8]),
	.C (op_a[5]),
	.B (op_a[7]),
	.A (op_a[6]) );
   NAND2X1 i_1041884 ( .Y (n_2088),
	.B (n_2017),
	.A (n_2087) );
   OAI211X1 i_834 ( .Y (n_2089),
	.C0 (cmd[1]),
	.B0 (op_b[9]),
	.A1 (cmd[0]),
	.A0 (op_a[9]) );
   OAI221XL i_836 ( .Y (n_2091),
	.C0 (n_2089),
	.B1 (n_3068),
	.B0 (n_1173),
	.A1 (n_1942),
	.A0 (n_1193) );
   AOI221X1 i_838 ( .Y (n_2093),
	.C0 (n_2091),
	.B1 (n_868),
	.B0 (n_1174),
	.A1 (op_a[9]),
	.A0 (n_2071) );
   OAI31X1 i_839 ( .Y (n_2094),
	.B0 (n_2093),
	.A2 (n_1264),
	.A1 (n_1738),
	.A0 (n_2079) );
   NAND2BX1 i_92 ( .Y (n_2096),
	.B (n_935),
	.AN (n_1776) );
   AOI21X1 i_1707216 ( .Y (n_2097),
	.B0 (n_1777),
	.A1 (n_1779),
	.A0 (n_1186) );
   NAND2X1 i_2027246 ( .Y (n_2098),
	.B (n_937),
	.A (n_1186) );
   OAI21XL i_1371491 ( .Y (n_2102),
	.B0 (n_1850),
	.A1 (n_1852),
	.A0 (n_1193) );
   NOR2X1 i_168 ( .Y (n_2103),
	.B (n_1147),
	.A (n_1193) );
   AOI21X1 i_93 ( .Y (n_2106),
	.B0 (n_1198),
	.A1 (op_b[10]),
	.A0 (op_a[10]) );
   NOR4BX1 i_1051885 ( .Y (n_2108),
	.D (n_2035),
	.C (op_a[9]),
	.B (op_a[8]),
	.AN (n_1887) );
   OAI211X1 i_866 ( .Y (n_2109),
	.C0 (cmd[1]),
	.B0 (op_b[10]),
	.A1 (cmd[0]),
	.A0 (op_a[10]) );
   OAI221XL i_868 ( .Y (n_2111),
	.C0 (n_2109),
	.B1 (n_3068),
	.B0 (n_1201),
	.A1 (n_1942),
	.A0 (n_1198) );
   AOI221X1 i_870 ( .Y (n_2113),
	.C0 (n_2111),
	.B1 (n_868),
	.B0 (n_1202),
	.A1 (op_a[10]),
	.A0 (n_2071) );
   OAI31X1 i_871 ( .Y (n_2114),
	.B0 (n_2113),
	.A2 (n_1287),
	.A1 (n_1738),
	.A0 (n_2096) );
   NAND2BX1 i_97 ( .Y (n_2116),
	.B (n_1237),
	.AN (n_1772) );
   AOI21X1 i_98 ( .Y (n_2118),
	.B0 (n_1244),
	.A1 (op_b[11]),
	.A0 (op_a[11]) );
   OAI211X1 i_896 ( .Y (n_2119),
	.C0 (cmd[1]),
	.B0 (op_b[11]),
	.A1 (cmd[0]),
	.A0 (op_a[11]) );
   OAI221XL i_898 ( .Y (n_2121),
	.C0 (n_2119),
	.B1 (n_3068),
	.B0 (n_1224),
	.A1 (n_1942),
	.A0 (n_1244) );
   AOI221X1 i_900 ( .Y (n_2123),
	.C0 (n_2121),
	.B1 (n_868),
	.B0 (n_1225),
	.A1 (op_a[11]),
	.A0 (n_2071) );
   OAI31X1 i_901 ( .Y (n_2124),
	.B0 (n_2123),
	.A2 (n_943),
	.A1 (n_1738),
	.A0 (n_2116) );
   NAND2BX1 i_102 ( .Y (n_2126),
	.B (n_933),
	.AN (n_1771) );
   AOI21X1 i_1727218 ( .Y (n_2127),
	.B0 (n_1772),
	.A1 (n_1776),
	.A0 (n_1237) );
   NAND2X1 i_2047248 ( .Y (n_2128),
	.B (n_935),
	.A (n_1237) );
   OAI21XL i_1391493 ( .Y (n_2132),
	.B0 (n_1845),
	.A1 (n_1849),
	.A0 (n_1244) );
   NOR2X1 i_170 ( .Y (n_2133),
	.B (n_1198),
	.A (n_1244) );
   AOI21X1 i_104 ( .Y (n_2136),
	.B0 (n_1249),
	.A1 (op_b[12]),
	.A0 (op_a[12]) );
   OAI211X1 i_928 ( .Y (n_2137),
	.C0 (cmd[1]),
	.B0 (op_b[12]),
	.A1 (cmd[0]),
	.A0 (op_a[12]) );
   OAI221XL i_930 ( .Y (n_2139),
	.C0 (n_2137),
	.B1 (n_3068),
	.B0 (n_1252),
	.A1 (n_1942),
	.A0 (n_1249) );
   AOI221X1 i_932 ( .Y (n_2141),
	.C0 (n_2139),
	.B1 (n_868),
	.B0 (n_1253),
	.A1 (op_a[12]),
	.A0 (n_2071) );
   OAI31X1 i_933 ( .Y (n_2142),
	.B0 (n_2141),
	.A2 (n_1334),
	.A1 (n_1738),
	.A0 (n_2126) );
   NAND2BX1 i_108 ( .Y (n_2144),
	.B (n_1286),
	.AN (n_1769) );
   AOI21X1 i_109 ( .Y (n_2150),
	.B0 (n_1293),
	.A1 (op_b[13]),
	.A0 (op_a[13]) );
   NOR4BX1 i_1081888 ( .Y (n_2153),
	.D (n_2088),
	.C (op_a[12]),
	.B (op_a[9]),
	.AN (n_1893) );
   OAI211X1 i_960 ( .Y (n_2154),
	.C0 (cmd[1]),
	.B0 (op_b[13]),
	.A1 (cmd[0]),
	.A0 (op_a[13]) );
   OAI221XL i_962 ( .Y (n_2156),
	.C0 (n_2154),
	.B1 (n_3068),
	.B0 (n_1273),
	.A1 (n_1942),
	.A0 (n_1293) );
   AOI221X1 i_964 ( .Y (n_2158),
	.C0 (n_2156),
	.B1 (n_868),
	.B0 (n_1274),
	.A1 (op_a[13]),
	.A0 (n_2071) );
   OAI31X1 i_965 ( .Y (n_2159),
	.B0 (n_2158),
	.A2 (n_1360),
	.A1 (n_1738),
	.A0 (n_2144) );
   NAND2BX1 i_113 ( .Y (n_2161),
	.B (n_931),
	.AN (n_1768) );
   AOI21X1 i_1747220 ( .Y (n_2162),
	.B0 (n_1769),
	.A1 (n_1771),
	.A0 (n_1286) );
   NAND2X1 i_2067250 ( .Y (n_2163),
	.B (n_933),
	.A (n_1286) );
   OAI21XL i_1411495 ( .Y (n_2167),
	.B0 (n_1842),
	.A1 (n_1844),
	.A0 (n_1293) );
   NOR2X1 i_172 ( .Y (n_2168),
	.B (n_1249),
	.A (n_1293) );
   AOI21X1 i_114 ( .Y (n_2171),
	.B0 (n_1297),
	.A1 (op_b[14]),
	.A0 (op_a[14]) );
   NOR4BBX1 i_1091889 ( .Y (n_2174),
	.D (op_a[13]),
	.C (op_a[12]),
	.BN (n_2108),
	.AN (n_1893) );
   OAI211X1 i_994 ( .Y (n_2175),
	.C0 (cmd[1]),
	.B0 (op_b[14]),
	.A1 (cmd[0]),
	.A0 (op_a[14]) );
   OAI221XL i_996 ( .Y (n_2177),
	.C0 (n_2175),
	.B1 (n_3068),
	.B0 (n_1300),
	.A1 (n_1942),
	.A0 (n_1297) );
   AOI221X1 i_998 ( .Y (n_2179),
	.C0 (n_2177),
	.B1 (n_868),
	.B0 (n_1301),
	.A1 (op_a[14]),
	.A0 (n_2071) );
   OAI31X1 i_999 ( .Y (n_2180),
	.B0 (n_2179),
	.A2 (n_1385),
	.A1 (n_1738),
	.A0 (n_2161) );
   NAND2BX1 i_118 ( .Y (n_2182),
	.B (n_1332),
	.AN (n_1764) );
   AOI21X1 i_119 ( .Y (n_2184),
	.B0 (n_1339),
	.A1 (op_b[15]),
	.A0 (op_a[15]) );
   OAI211X1 i_1018 ( .Y (n_2185),
	.C0 (cmd[1]),
	.B0 (op_b[15]),
	.A1 (cmd[0]),
	.A0 (op_a[15]) );
   OAI221XL i_1020 ( .Y (n_2187),
	.C0 (n_2185),
	.B1 (n_3068),
	.B0 (n_1319),
	.A1 (n_1942),
	.A0 (n_1339) );
   AOI221X1 i_1022 ( .Y (n_2189),
	.C0 (n_2187),
	.B1 (n_868),
	.B0 (n_1320),
	.A1 (op_a[15]),
	.A0 (n_2071) );
   OAI31X1 i_1023 ( .Y (n_2190),
	.B0 (n_2189),
	.A2 (n_1411),
	.A1 (n_1738),
	.A0 (n_2182) );
   NAND2BX1 i_123 ( .Y (n_2192),
	.B (n_929),
	.AN (n_1763) );
   AOI21X1 i_1767222 ( .Y (n_2193),
	.B0 (n_1764),
	.A1 (n_1768),
	.A0 (n_1332) );
   NAND2X1 i_2087252 ( .Y (n_2194),
	.B (n_931),
	.A (n_1332) );
   OAI21XL i_1431497 ( .Y (n_2198),
	.B0 (n_1837),
	.A1 (n_1841),
	.A0 (n_1339) );
   NOR2X1 i_174 ( .Y (n_2199),
	.B (n_1297),
	.A (n_1339) );
   AOI21X1 i_124 ( .Y (n_2202),
	.B0 (n_1344),
	.A1 (op_b[16]),
	.A0 (op_a[16]) );
   OAI211X1 i_1051 ( .Y (n_2203),
	.C0 (cmd[1]),
	.B0 (op_b[16]),
	.A1 (cmd[0]),
	.A0 (op_a[16]) );
   OAI221XL i_1053 ( .Y (n_2205),
	.C0 (n_2203),
	.B1 (n_3068),
	.B0 (n_1347),
	.A1 (n_1942),
	.A0 (n_1344) );
   AOI221X1 i_1055 ( .Y (n_2207),
	.C0 (n_2205),
	.B1 (n_868),
	.B0 (n_1348),
	.A1 (op_a[16]),
	.A0 (n_2071) );
   OAI31X1 i_1056 ( .Y (n_2208),
	.B0 (n_2207),
	.A2 (n_1436),
	.A1 (n_1738),
	.A0 (n_2192) );
   NAND2BX1 i_128 ( .Y (n_2210),
	.B (n_1383),
	.AN (n_1761) );
   AOI21X1 i_129 ( .Y (n_2216),
	.B0 (n_1390),
	.A1 (op_b[17]),
	.A0 (op_a[17]) );
   NOR4X1 i_1067 ( .Y (n_2218),
	.D (op_a[16]),
	.C (op_a[15]),
	.B (op_a[14]),
	.A (op_a[13]) );
   NAND2X1 i_1441918 ( .Y (n_2219),
	.B (n_2153),
	.A (n_2218) );
   OAI211X1 i_1089 ( .Y (n_2220),
	.C0 (cmd[1]),
	.B0 (op_b[17]),
	.A1 (cmd[0]),
	.A0 (op_a[17]) );
   OAI221XL i_1091 ( .Y (n_2222),
	.C0 (n_2220),
	.B1 (n_3068),
	.B0 (n_1370),
	.A1 (n_1942),
	.A0 (n_1390) );
   AOI221X1 i_1094 ( .Y (n_2224),
	.C0 (n_2222),
	.B1 (n_868),
	.B0 (n_1371),
	.A1 (op_a[17]),
	.A0 (n_2071) );
   OAI31X1 i_1096 ( .Y (n_2225),
	.B0 (n_2224),
	.A2 (n_1462),
	.A1 (n_1738),
	.A0 (n_2210) );
   NAND2BX1 i_133 ( .Y (n_2227),
	.B (n_927),
	.AN (n_1760) );
   AOI21X1 i_1787224 ( .Y (n_2228),
	.B0 (n_1761),
	.A1 (n_1763),
	.A0 (n_1383) );
   NAND2X1 i_2107254 ( .Y (n_2229),
	.B (n_929),
	.A (n_1383) );
   OAI21XL i_1451499 ( .Y (n_2233),
	.B0 (n_1834),
	.A1 (n_1836),
	.A0 (n_1390) );
   NOR2X1 i_176 ( .Y (n_2234),
	.B (n_1344),
	.A (n_1390) );
   AOI21X1 i_134 ( .Y (n_2237),
	.B0 (n_1395),
	.A1 (op_b[18]),
	.A0 (op_a[18]) );
   NOR4X1 i_1111 ( .Y (n_2239),
	.D (op_a[15]),
	.C (op_a[14]),
	.B (op_a[17]),
	.A (op_a[16]) );
   OAI211X1 i_1132 ( .Y (n_2241),
	.C0 (cmd[1]),
	.B0 (op_b[18]),
	.A1 (cmd[0]),
	.A0 (op_a[18]) );
   OAI221XL i_1134 ( .Y (n_2243),
	.C0 (n_2241),
	.B1 (n_3068),
	.B0 (n_1398),
	.A1 (n_1942),
	.A0 (n_1395) );
   AOI221X1 i_1137 ( .Y (n_2245),
	.C0 (n_2243),
	.B1 (n_868),
	.B0 (n_1399),
	.A1 (op_a[18]),
	.A0 (n_2071) );
   OAI31X1 i_1138 ( .Y (n_2246),
	.B0 (n_2245),
	.A2 (n_1487),
	.A1 (n_1738),
	.A0 (n_2227) );
   NAND2BX1 i_190 ( .Y (n_2248),
	.B (n_1434),
	.AN (n_1756) );
   AOI21X1 i_191 ( .Y (n_2250),
	.B0 (n_1441),
	.A1 (op_b[19]),
	.A0 (op_a[19]) );
   OAI211X1 i_1168 ( .Y (n_2251),
	.C0 (cmd[1]),
	.B0 (op_b[19]),
	.A1 (cmd[0]),
	.A0 (op_a[19]) );
   OAI221XL i_1170 ( .Y (n_2253),
	.C0 (n_2251),
	.B1 (n_3068),
	.B0 (n_1421),
	.A1 (n_1942),
	.A0 (n_1441) );
   AOI221X1 i_1173 ( .Y (n_2255),
	.C0 (n_2253),
	.B1 (n_868),
	.B0 (n_1422),
	.A1 (op_a[19]),
	.A0 (n_2071) );
   OAI31X1 i_1174 ( .Y (n_2256),
	.B0 (n_2255),
	.A2 (n_946),
	.A1 (n_1738),
	.A0 (n_2248) );
   NAND2BX1 i_222 ( .Y (n_2258),
	.B (n_925),
	.AN (n_1755) );
   AOI21X1 i_1807226 ( .Y (n_2259),
	.B0 (n_1756),
	.A1 (n_1760),
	.A0 (n_1434) );
   NAND2X1 i_2127256 ( .Y (n_2260),
	.B (n_927),
	.A (n_1434) );
   OAI21XL i_1471501 ( .Y (n_2264),
	.B0 (n_1829),
	.A1 (n_1833),
	.A0 (n_1441) );
   NOR2X1 i_178 ( .Y (n_2265),
	.B (n_1395),
	.A (n_1441) );
   AOI21X1 i_224 ( .Y (n_2268),
	.B0 (n_1446),
	.A1 (op_b[20]),
	.A0 (op_a[20]) );
   OAI211X1 i_1206 ( .Y (n_2269),
	.C0 (cmd[1]),
	.B0 (op_b[20]),
	.A1 (cmd[0]),
	.A0 (op_a[20]) );
   OAI221XL i_1209 ( .Y (n_2271),
	.C0 (n_2269),
	.B1 (n_3068),
	.B0 (n_1449),
	.A1 (n_1942),
	.A0 (n_1446) );
   AOI221X1 i_1211 ( .Y (n_2273),
	.C0 (n_2271),
	.B1 (n_868),
	.B0 (n_1450),
	.A1 (op_a[20]),
	.A0 (n_2071) );
   OAI31X1 i_1212 ( .Y (n_2274),
	.B0 (n_2273),
	.A2 (n_1534),
	.A1 (n_1738),
	.A0 (n_2258) );
   NAND2BX1 i_229 ( .Y (n_2276),
	.B (n_1485),
	.AN (n_1753) );
   AOI21X1 i_230 ( .Y (n_2282),
	.B0 (n_1492),
	.A1 (op_b[21]),
	.A0 (op_a[21]) );
   NOR4BX1 i_1481922 ( .Y (n_2285),
	.D (n_2219),
	.C (op_a[20]),
	.B (op_a[17]),
	.AN (n_1901) );
   OAI211X1 i_1245 ( .Y (n_2286),
	.C0 (cmd[1]),
	.B0 (op_b[21]),
	.A1 (cmd[0]),
	.A0 (op_a[21]) );
   OAI221XL i_1247 ( .Y (n_2288),
	.C0 (n_2286),
	.B1 (n_3068),
	.B0 (n_1472),
	.A1 (n_1942),
	.A0 (n_1492) );
   AOI221X1 i_1249 ( .Y (n_2290),
	.C0 (n_2288),
	.B1 (n_868),
	.B0 (n_1473),
	.A1 (op_a[21]),
	.A0 (n_2071) );
   OAI31X1 i_1250 ( .Y (n_2291),
	.B0 (n_2290),
	.A2 (n_1561),
	.A1 (n_1738),
	.A0 (n_2276) );
   NAND2BX1 i_236 ( .Y (n_2293),
	.B (n_923),
	.AN (n_1752) );
   AOI21X1 i_1827228 ( .Y (n_2294),
	.B0 (n_1753),
	.A1 (n_1755),
	.A0 (n_1485) );
   NAND2X1 i_2147258 ( .Y (n_2295),
	.B (n_925),
	.A (n_1485) );
   OAI21XL i_1491503 ( .Y (n_2299),
	.B0 (n_1826),
	.A1 (n_1828),
	.A0 (n_1492) );
   NOR2X1 i_180 ( .Y (n_2300),
	.B (n_1446),
	.A (n_1492) );
   AOI21X1 i_237 ( .Y (n_2303),
	.B0 (n_1497),
	.A1 (op_b[22]),
	.A0 (op_a[22]) );
   NAND4X1 i_1491923 ( .Y (n_2305),
	.D (n_2174),
	.C (n_2239),
	.B (n_1901),
	.A (n_1905) );
   OAI211X1 i_1284 ( .Y (n_2306),
	.C0 (cmd[1]),
	.B0 (op_b[22]),
	.A1 (cmd[0]),
	.A0 (op_a[22]) );
   OAI221XL i_1286 ( .Y (n_2308),
	.C0 (n_2306),
	.B1 (n_3068),
	.B0 (n_1500),
	.A1 (n_1942),
	.A0 (n_1497) );
   AOI221X1 i_1289 ( .Y (n_2310),
	.C0 (n_2308),
	.B1 (n_868),
	.B0 (n_1501),
	.A1 (op_a[22]),
	.A0 (n_2071) );
   OAI31X1 i_1290 ( .Y (n_2311),
	.B0 (n_2310),
	.A2 (n_1587),
	.A1 (n_1738),
	.A0 (n_2293) );
   NAND2BX1 i_242 ( .Y (n_2313),
	.B (n_1532),
	.AN (n_1748) );
   AOI21X1 i_244 ( .Y (n_2315),
	.B0 (n_1539),
	.A1 (op_b[23]),
	.A0 (op_a[23]) );
   OAI211X1 i_1311 ( .Y (n_2316),
	.C0 (cmd[1]),
	.B0 (op_b[23]),
	.A1 (cmd[0]),
	.A0 (op_a[23]) );
   OAI221XL i_1313 ( .Y (n_2318),
	.C0 (n_2316),
	.B1 (n_3068),
	.B0 (n_1519),
	.A1 (n_1942),
	.A0 (n_1539) );
   AOI221X1 i_1316 ( .Y (n_2320),
	.C0 (n_2318),
	.B1 (n_868),
	.B0 (n_1520),
	.A1 (op_a[23]),
	.A0 (n_2071) );
   OAI31X1 i_1317 ( .Y (n_2321),
	.B0 (n_2320),
	.A2 (n_1612),
	.A1 (n_1738),
	.A0 (n_2313) );
   NAND2BX1 i_249 ( .Y (n_2323),
	.B (n_921),
	.AN (n_1747) );
   AOI21X1 i_1847230 ( .Y (n_2324),
	.B0 (n_1748),
	.A1 (n_1752),
	.A0 (n_1532) );
   NAND2X1 i_2167260 ( .Y (n_2325),
	.B (n_923),
	.A (n_1532) );
   OAI21XL i_1511505 ( .Y (n_2329),
	.B0 (n_1821),
	.A1 (n_1825),
	.A0 (n_1539) );
   NOR2X1 i_182 ( .Y (n_2330),
	.B (n_1497),
	.A (n_1539) );
   AOI21X1 i_250 ( .Y (n_2333),
	.B0 (n_1544),
	.A1 (op_b[24]),
	.A0 (op_a[24]) );
   OAI211X1 i_1349 ( .Y (n_2334),
	.C0 (cmd[1]),
	.B0 (op_b[24]),
	.A1 (cmd[0]),
	.A0 (op_a[24]) );
   OAI221XL i_1352 ( .Y (n_2336),
	.C0 (n_2334),
	.B1 (n_3068),
	.B0 (n_1547),
	.A1 (n_1942),
	.A0 (n_1544) );
   AOI221X1 i_1354 ( .Y (n_2338),
	.C0 (n_2336),
	.B1 (n_868),
	.B0 (n_1548),
	.A1 (op_a[24]),
	.A0 (n_2071) );
   OAI31X1 i_1355 ( .Y (n_2339),
	.B0 (n_2338),
	.A2 (n_1637),
	.A1 (n_1738),
	.A0 (n_2323) );
   NAND2BX1 i_255 ( .Y (n_2341),
	.B (n_1585),
	.AN (n_1745) );
   OAI21XL i_2487288 ( .Y (n_2342),
	.B0 (n_1749),
	.A1 (n_1808),
	.A0 (n_1754) );
   AOI31X1 i_4377415 ( .Y (n_2344),
	.B0 (n_2342),
	.A2 (n_1758),
	.A1 (n_3071),
	.A0 (n_1561) );
   AOI21X1 i_214 ( .Y (n_2346),
	.B0 (n_1822),
	.A1 (n_1881),
	.A0 (n_1827) );
   AOI21X1 i_260 ( .Y (n_2349),
	.B0 (n_1592),
	.A1 (op_b[25]),
	.A0 (op_a[25]) );
   NOR4X1 i_1367 ( .Y (n_2351),
	.D (op_a[24]),
	.C (op_a[21]),
	.B (op_a[23]),
	.A (op_a[22]) );
   NAND2X1 i_1521926 ( .Y (n_2352),
	.B (n_2285),
	.A (n_2351) );
   OAI211X1 i_1399 ( .Y (n_2353),
	.C0 (cmd[1]),
	.B0 (op_b[25]),
	.A1 (cmd[0]),
	.A0 (op_a[25]) );
   OAI221XL i_1401 ( .Y (n_2355),
	.C0 (n_2353),
	.B1 (n_3068),
	.B0 (n_1572),
	.A1 (n_1942),
	.A0 (n_1592) );
   AOI211X1 i_1403 ( .Y (n_2357),
	.C0 (n_1579),
	.B0 (n_2355),
	.A1 (op_a[25]),
	.A0 (n_2071) );
   OAI31X1 i_1404 ( .Y (n_2358),
	.B0 (n_2357),
	.A2 (n_1738),
	.A1 (n_2341),
	.A0 (n_3093) );
   NAND2BX1 i_264 ( .Y (n_2360),
	.B (n_1709),
	.AN (n_1744) );
   AOI21X1 i_1867232 ( .Y (n_2361),
	.B0 (n_1745),
	.A1 (n_1747),
	.A0 (n_1585) );
   AND2X1 i_2187262 ( .Y (n_2362),
	.B (n_921),
	.A (n_1585) );
   OAI21XL i_1531507 ( .Y (n_2366),
	.B0 (n_1818),
	.A1 (n_1820),
	.A0 (n_1592) );
   NOR2X1 i_184 ( .Y (n_2367),
	.B (n_1544),
	.A (n_1592) );
   AOI21X1 i_265 ( .Y (n_2370),
	.B0 (n_1700),
	.A1 (op_b[26]),
	.A0 (op_a[26]) );
   NOR4BX1 i_1531927 ( .Y (n_2372),
	.D (n_2305),
	.C (op_a[25]),
	.B (op_a[24]),
	.AN (n_1904) );
   OAI211X1 i_1435 ( .Y (n_2373),
	.C0 (cmd[1]),
	.B0 (op_b[26]),
	.A1 (cmd[0]),
	.A0 (op_a[26]) );
   OAI221XL i_1437 ( .Y (n_2375),
	.C0 (n_2373),
	.B1 (n_3068),
	.B0 (n_1599),
	.A1 (n_1942),
	.A0 (n_1700) );
   AOI221X1 i_1439 ( .Y (n_2377),
	.C0 (n_2375),
	.B1 (n_868),
	.B0 (n_1600),
	.A1 (op_a[26]),
	.A0 (n_2071) );
   OAI31X1 i_1440 ( .Y (n_2378),
	.B0 (n_2377),
	.A2 (n_1708),
	.A1 (n_1738),
	.A0 (n_2360) );
   AOI21X1 i_271 ( .Y (n_2382),
	.B0 (n_1650),
	.A1 (op_b[27]),
	.A0 (op_a[27]) );
   OAI211X1 i_1465 ( .Y (n_2383),
	.C0 (cmd[1]),
	.B0 (op_b[27]),
	.A1 (cmd[0]),
	.A0 (op_a[27]) );
   OAI21XL i_1466 ( .Y (n_2384),
	.B0 (n_2383),
	.A1 (n_1942),
	.A0 (n_1650) );
   AOI21X1 i_1467 ( .Y (n_2385),
	.B0 (n_2384),
	.A1 (op_a[27]),
	.A0 (n_2071) );
   OAI221XL i_1469 ( .Y (n_2387),
	.C0 (n_2385),
	.B1 (n_3095),
	.B0 (n_1623),
	.A1 (n_1622),
	.A0 (n_3068) );
   NOR2BX1 i_276 ( .Y (n_2390),
	.B (n_1710),
	.AN (n_1706) );
   OAI2BB1X1 i_1887234 ( .Y (n_2391),
	.B0 (n_3069),
	.A1N (n_1744),
	.A0N (n_1640) );
   AOI31X1 i_440 ( .Y (n_2393),
	.B0 (n_2391),
	.A2 (n_1639),
	.A1 (n_1709),
	.A0 (n_1640) );
   OAI211X1 i_1501 ( .Y (n_2394),
	.C0 (cmd[1]),
	.B0 (op_b[28]),
	.A1 (cmd[0]),
	.A0 (op_a[28]) );
   OAI2BB1X1 i_1502 ( .Y (n_2395),
	.B0 (n_2394),
	.A1N (n_3064),
	.A0N (n_3066) );
   AOI211X1 i_1504 ( .Y (n_2397),
	.C0 (n_1661),
	.B0 (n_2395),
	.A1 (op_a[28]),
	.A0 (n_2071) );
   OAI21XL i_1551509 ( .Y (n_2399),
	.B0 (n_1814),
	.A1 (n_1817),
	.A0 (n_1650) );
   NOR2BX1 i_403 ( .Y (n_2401),
	.B (n_2399),
	.AN (n_1648) );
   AOI21X1 i_277 ( .Y (n_2402),
	.B0 (n_1697),
	.A1 (op_b[28]),
	.A0 (op_a[28]) );
   AOI32X1 i_1506 ( .Y (n_2404),
	.B1 (n_868),
	.B0 (n_1656),
	.A2 (n_2390),
	.A1 (n_3062),
	.A0 (n_2393) );
   NAND2BX1 i_281 ( .Y (n_2406),
	.B (n_885),
	.AN (n_1713) );
   OAI21XL i_1514 ( .Y (n_2408),
	.B0 (n_1746),
	.A1 (n_3090),
	.A0 (n_1750) );
   OAI21XL i_441 ( .Y (n_2409),
	.B0 (n_1742),
	.A1 (n_1743),
	.A0 (n_1670) );
   AOI21X1 i_1524 ( .Y (n_2411),
	.B0 (n_1819),
	.A1 (n_3091),
	.A0 (n_1823) );
   OAI21XL i_283 ( .Y (n_2413),
	.B0 (n_1812),
	.A1 (op_a[29]),
	.A0 (op_b[29]) );
   NOR4BX1 i_1561930 ( .Y (n_2417),
	.D (n_2352),
	.C (op_a[28]),
	.B (op_a[25]),
	.AN (n_1908) );
   OAI211X1 i_1537 ( .Y (n_2418),
	.C0 (cmd[1]),
	.B0 (op_b[29]),
	.A1 (cmd[0]),
	.A0 (op_a[29]) );
   OAI221XL i_1539 ( .Y (n_2420),
	.C0 (n_2418),
	.B1 (n_3068),
	.B0 (n_1682),
	.A1 (n_1942),
	.A0 (n_1703) );
   AOI211X1 i_1541 ( .Y (n_2422),
	.C0 (n_1689),
	.B0 (n_2420),
	.A1 (op_a[29]),
	.A0 (n_2071) );
   OAI2BB1X1 i_1542 ( .Y (n_2423),
	.B0 (n_2422),
	.A1N (n_868),
	.A0N (n_1683) );
   NAND2BX1 i_1587204 ( .Y (n_2425),
	.B (n_954),
	.AN (n_952) );
   NOR2BX1 i_1565 ( .Y (n_2426),
	.B (n_1743),
	.AN (n_1709) );
   OAI21XL i_442 ( .Y (n_2428),
	.B0 (n_885),
	.A1 (n_1713),
	.A0 (n_1714) );
   OAI21XL i_405 ( .Y (n_2431),
	.B0 (n_1812),
	.A1 (n_1703),
	.A0 (n_1704) );
   NAND3X1 i_1571931 ( .Y (n_2434),
	.C (n_2372),
	.B (n_1908),
	.A (n_1912) );
   AOI211X1 i_1553 ( .Y (n_2436),
	.C0 (n_3064),
	.B0 (n_2071),
	.A1 (op_b[30]),
	.A0 (cmd[1]) );
   NOR2BX1 i_1578 ( .Y (n_2437),
	.B (op_a[30]),
	.AN (n_2434) );
   AOI222X1 i_1580 ( .Y (n_2439),
	.C1 (op_a[30]),
	.C0 (n_1720),
	.B1 (n_1946),
	.B0 (op_b[30]),
	.A1 (n_1918),
	.A0 (n_2437) );
   OAI221XL i_1582 ( .Y (n_2441),
	.C0 (n_2439),
	.B1 (n_2425),
	.B0 (n_1723),
	.A1 (n_3068),
	.A0 (n_1915) );
   NOR4X1 i_81615 ( .Y (n_868),
	.D (cmd[1]),
	.C (cmd[3]),
	.B (cmd[2]),
	.A (cmd[0]) );
   AOI21X1 i_1398 ( .Y (result[32]),
	.B0 (n_828),
	.A1 (n_3095),
	.A0 (n_1738) );
   NOR4BBX1 i_671598 ( .Y (n_166),
	.D (n_1911),
	.C (op_a[30]),
	.BN (op_a[31]),
	.AN (n_1912) );
   NAND2X1 i_2154 ( .Y (n_9076575),
	.B (result[32]),
	.A (ovm) );
   INVX1 i_3032 ( .Y (n_3060),
	.A (n_827) );
   INVX1 i_3034 ( .Y (n_3062),
	.A (n_1738) );
   INVX1 i_3035 ( .Y (n_3063),
	.A (n_1944) );
   INVX1 i_3036 ( .Y (n_3064),
	.A (n_1942) );
   INVX1 i_3037 ( .Y (n_3065),
	.A (n_1136) );
   INVX1 i_3038 ( .Y (n_3066),
	.A (n_1697) );
   INVX1 i_3039 ( .Y (n_3067),
	.A (n_1886) );
   INVX1 i_3040 ( .Y (n_3068),
	.A (n_1918) );
   INVX1 i_3041 ( .Y (n_3069),
	.A (n_1741) );
   INVX1 i_3042 ( .Y (n_3070),
	.A (n_1742) );
   INVX1 i_3043 ( .Y (n_3071),
	.A (n_1808) );
   INVX1 i_3044 ( .Y (result[0]),
	.A (n_984) );
   INVX1 i_3045 ( .Y (n_3073),
	.A (n_1781) );
   INVX1 i_3046 ( .Y (n_3074),
	.A (n_1784) );
   INVX1 i_3047 ( .Y (n_3075),
	.A (n_1793) );
   INVX1 i_3048 ( .Y (n_3076),
	.A (n_1213) );
   INVX1 i_3049 ( .Y (n_3077),
	.A (n_1816) );
   INVX1 i_3050 ( .Y (n_3078),
	.A (n_1853) );
   INVX1 i_3051 ( .Y (n_3079),
	.A (n_1858) );
   INVX1 i_3052 ( .Y (n_3080),
	.A (n_1857) );
   INVX1 i_3053 ( .Y (n_3081),
	.A (n_1861) );
   INVX1 i_3054 ( .Y (n_3082),
	.A (n_1860) );
   INVX1 i_3055 ( .Y (n_3083),
	.A (n_1866) );
   INVX1 i_3056 ( .Y (n_3084),
	.A (n_1865) );
   INVX1 i_3057 ( .Y (n_3085),
	.A (n_1868) );
   INVX1 i_3058 ( .Y (n_3086),
	.A (n_911) );
   INVX1 i_3059 ( .Y (n_3087),
	.A (n_1996) );
   INVX1 i_3060 ( .Y (n_3088),
	.A (n_2428) );
   INVX1 i_3061 ( .Y (n_3089),
	.A (n_2040) );
   INVX1 i_3062 ( .Y (n_3090),
	.A (n_2342) );
   INVX1 i_3063 ( .Y (n_3091),
	.A (n_2346) );
   INVX1 i_3064 ( .Y (n_3092),
	.A (n_2083) );
   INVX1 i_3065 ( .Y (n_3093),
	.A (n_2344) );
   INVX1 i_3066 ( .Y (n_907),
	.A (n_9076575) );
   INVX1 i_3067 ( .Y (n_3095),
	.A (n_868) );
endmodule

module data_bus_mach (
	clk,
	reset,
	read,
	write,
	address,
	data_in,
	data_out,
	pad_data_in,
	pad_data_out,
	addrs_in,
	read_cycle,
	sync,
	go,
	as,
	done,
	bus_request,
	bus_grant,
	scan_en,
	BG_scan_in,
	BG_scan_out );
   input clk;
   input reset;
   output read;
   output write;
   output [7:0] address;
   input [15:0] data_in;
   output [15:0] data_out;
   input [15:0] pad_data_in;
   output [15:0] pad_data_out;
   input [7:0] addrs_in;
   input read_cycle;
   input sync;
   input go;
   output as;
   output done;
   output bus_request;
   input bus_grant;
   input scan_en;
   input BG_scan_in;
   output BG_scan_out;

   // Internal wires
   wire [2:0] present_state;
   wire n_7893;
   wire n_6389;
   wire FE_OFN88_tdsp_data_out_0_;
   wire FE_OFN84_tdsp_data_out_1_;
   wire n_6381;
   wire FE_OFN81_tdsp_data_out_2_;
   wire FE_OFN76_tdsp_data_out_3_;
   wire n_6373;
   wire FE_OFN71_tdsp_data_out_4_;
   wire FE_OFN66_tdsp_data_out_5_;
   wire FE_OFN62_tdsp_data_out_6_;
   wire n_6361;
   wire FE_OFN53_tdsp_data_out_8_;
   wire FE_OFN48_tdsp_data_out_9_;
   wire n_6353;
   wire FE_OFN44_tdsp_data_out_10_;
   wire n_6349;
   wire FE_OFN40_tdsp_data_out_11_;
   wire FE_OFN35_tdsp_data_out_12_;
   wire n_6341;
   wire FE_OFN30_tdsp_data_out_13_;
   wire n_6337;
   wire FE_OFN25_tdsp_data_out_14_;
   wire n_6333;
   wire FE_OFN22_tdsp_data_out_15_;
   wire n_6329;
   wire FE_OFN107_t_addrs_1_;
   wire n_6325;
   wire n_6321;
   wire n_6317;
   wire n_6313;
   wire FE_OFN110_t_addrs_0_;
   wire FE_OFN101_t_addrs_3_;
   wire FE_OFN104_t_addrs_2_;
   wire FE_OFN57_tdsp_data_out_7_;
   wire n_16;
   wire n_23;
   wire n_21;
   wire \nbus_626[0] ;
   wire n_4642;
   wire FE_OFN6_scan_enI;
   wire n_4641;
   wire n_24;
   wire n_4534;
   wire n_5177;
   wire n_4540;
   wire n_4546;
   wire n_28;
   wire n_5205;
   wire n_4640;
   wire n_4552;
   wire n_4558;
   wire n_4564;
   wire n_4570;
   wire n_4576;
   wire FE_OFN135_scan_enI;
   wire n_4582;
   wire FE_OFN19_scan_enI;
   wire n_4588;
   wire n_31;
   wire n_4594;
   wire n_4600;
   wire n_5232;
   wire n_4606;
   wire n_5226;
   wire n_4612;
   wire n_4618;
   wire n_4624;
   wire FE_OFN149_tdsp_data_out_15_;
   wire FE_OFN111_t_addrs_0_;
   wire FE_OFN108_t_addrs_1_;
   wire FE_OFN105_t_addrs_2_;
   wire FE_OFN102_t_addrs_3_;
   wire FE_OFN77_tdsp_data_out_3_;
   wire FE_OFN72_tdsp_data_out_4_;
   wire FE_OFN67_tdsp_data_out_5_;
   wire FE_OFN54_tdsp_data_out_8_;
   wire FE_OFN36_tdsp_data_out_12_;
   wire FE_OFN31_tdsp_data_out_13_;

   INVXL i_10642 ( .Y (BG_scan_out),
	.A (n_7893) );
   INVXL i_10641 ( .Y (n_7893),
	.A (bus_request) );
   INVXL i_9590 ( .Y (FE_OFN88_tdsp_data_out_0_),
	.A (n_6389) );
   INVXL i_9589 ( .Y (n_6389),
	.A (data_in[0]) );
   BUFX3 i_9588 ( .Y (FE_OFN84_tdsp_data_out_1_),
	.A (data_in[1]) );
   INVXL i_9584 ( .Y (FE_OFN81_tdsp_data_out_2_),
	.A (n_6381) );
   INVXL i_9583 ( .Y (n_6381),
	.A (data_in[2]) );
   CLKBUFX2 i_9582 ( .Y (FE_OFN76_tdsp_data_out_3_),
	.A (data_in[3]) );
   INVXL i_9578 ( .Y (FE_OFN71_tdsp_data_out_4_),
	.A (n_6373) );
   INVXL i_9577 ( .Y (n_6373),
	.A (data_in[4]) );
   BUFX3 i_9576 ( .Y (FE_OFN66_tdsp_data_out_5_),
	.A (data_in[5]) );
   BUFX3 i_9573 ( .Y (FE_OFN62_tdsp_data_out_6_),
	.A (data_in[6]) );
   INVX1 i_9569 ( .Y (FE_OFN53_tdsp_data_out_8_),
	.A (n_6361) );
   INVXL i_9568 ( .Y (n_6361),
	.A (data_in[8]) );
   BUFX3 i_9567 ( .Y (FE_OFN48_tdsp_data_out_9_),
	.A (data_in[9]) );
   INVXL i_9563 ( .Y (FE_OFN44_tdsp_data_out_10_),
	.A (n_6353) );
   INVXL i_9562 ( .Y (n_6353),
	.A (data_in[10]) );
   INVXL i_9560 ( .Y (FE_OFN40_tdsp_data_out_11_),
	.A (n_6349) );
   INVXL i_9559 ( .Y (n_6349),
	.A (data_in[11]) );
   CLKBUFX2 i_9558 ( .Y (FE_OFN35_tdsp_data_out_12_),
	.A (data_in[12]) );
   INVXL i_9554 ( .Y (FE_OFN30_tdsp_data_out_13_),
	.A (n_6341) );
   INVXL i_9553 ( .Y (n_6341),
	.A (data_in[13]) );
   INVX1 i_9551 ( .Y (FE_OFN25_tdsp_data_out_14_),
	.A (n_6337) );
   INVXL i_9550 ( .Y (n_6337),
	.A (data_in[14]) );
   INVX2 i_9548 ( .Y (FE_OFN22_tdsp_data_out_15_),
	.A (n_6333) );
   INVXL i_9547 ( .Y (n_6333),
	.A (data_in[15]) );
   INVXL i_9545 ( .Y (FE_OFN107_t_addrs_1_),
	.A (n_6329) );
   INVXL i_9544 ( .Y (n_6329),
	.A (addrs_in[1]) );
   INVX2 i_9542 ( .Y (address[4]),
	.A (n_6325) );
   INVXL i_9541 ( .Y (n_6325),
	.A (addrs_in[4]) );
   INVX2 i_9539 ( .Y (address[5]),
	.A (n_6321) );
   INVXL i_9538 ( .Y (n_6321),
	.A (addrs_in[5]) );
   INVX2 i_9536 ( .Y (address[6]),
	.A (n_6317) );
   INVXL i_9535 ( .Y (n_6317),
	.A (addrs_in[6]) );
   INVXL i_9533 ( .Y (address[7]),
	.A (n_6313) );
   INVXL i_9532 ( .Y (n_6313),
	.A (addrs_in[7]) );
   CLKBUFX1 i_9491 ( .Y (FE_OFN110_t_addrs_0_),
	.A (addrs_in[0]) );
   CLKBUFX2 i_9486 ( .Y (FE_OFN101_t_addrs_3_),
	.A (addrs_in[3]) );
   CLKBUFX2 i_9485 ( .Y (FE_OFN104_t_addrs_2_),
	.A (addrs_in[2]) );
   CLKBUFX2 i_9474 ( .Y (FE_OFN57_tdsp_data_out_7_),
	.A (data_in[7]) );
   NOR2X1 i_11 ( .Y (n_16),
	.B (present_state[2]),
	.A (go) );
   OAI21XL i_8 ( .Y (n_21),
	.B0 (n_23),
	.A1 (present_state[1]),
	.A0 (n_16) );
   SDFFRHQX1 present_state_reg_0 ( .SI (BG_scan_in),
	.SE (scan_en),
	.RN (n_4642),
	.Q (present_state[0]),
	.D (\nbus_626[0] ),
	.CK (clk) );
   SDFFRHQX1 present_state_reg_1 ( .SI (present_state[0]),
	.SE (FE_OFN6_scan_enI),
	.RN (n_4642),
	.Q (present_state[1]),
	.D (n_4641),
	.CK (clk) );
   SDFFRHQX1 present_state_reg_2 ( .SI (present_state[1]),
	.SE (scan_en),
	.RN (n_4642),
	.Q (present_state[2]),
	.D (n_24),
	.CK (clk) );
   SDFFRHQX1 data_out_reg_0 ( .SI (present_state[2]),
	.SE (scan_en),
	.RN (n_4642),
	.Q (data_out[0]),
	.D (n_4534),
	.CK (clk) );
   MX2X1 i_6145 ( .Y (n_4534),
	.S0 (n_5177),
	.B (pad_data_in[0]),
	.A (data_out[0]) );
   SDFFRHQX1 data_out_reg_1 ( .SI (data_out[0]),
	.SE (scan_en),
	.RN (n_4642),
	.Q (data_out[1]),
	.D (n_4540),
	.CK (clk) );
   MX2X1 i_6152 ( .Y (n_4540),
	.S0 (n_5177),
	.B (pad_data_in[1]),
	.A (data_out[1]) );
   XNOR2X1 i_3 ( .Y (n_23),
	.B (present_state[1]),
	.A (present_state[0]) );
   SDFFRHQX1 data_out_reg_2 ( .SI (data_out[1]),
	.SE (scan_en),
	.RN (n_4642),
	.Q (data_out[2]),
	.D (n_4546),
	.CK (clk) );
   MX2X1 i_6159 ( .Y (n_4546),
	.S0 (n_5177),
	.B (pad_data_in[2]),
	.A (data_out[2]) );
   OAI32X1 i_2 ( .Y (n_24),
	.B1 (n_4640),
	.B0 (n_5205),
	.A2 (n_28),
	.A1 (present_state[0]),
	.A0 (present_state[1]) );
   SDFFRHQX1 data_out_reg_3 ( .SI (data_out[2]),
	.SE (scan_en),
	.RN (n_4642),
	.Q (data_out[3]),
	.D (n_4552),
	.CK (clk) );
   MX2X1 i_6166 ( .Y (n_4552),
	.S0 (n_5177),
	.B (pad_data_in[3]),
	.A (data_out[3]) );
   SDFFRHQX1 data_out_reg_4 ( .SI (data_out[3]),
	.SE (scan_en),
	.RN (n_4642),
	.Q (data_out[4]),
	.D (n_4558),
	.CK (clk) );
   MX2X1 i_6173 ( .Y (n_4558),
	.S0 (n_5177),
	.B (pad_data_in[4]),
	.A (data_out[4]) );
   SDFFRHQX1 data_out_reg_5 ( .SI (data_out[4]),
	.SE (FE_OFN6_scan_enI),
	.RN (n_4642),
	.Q (data_out[5]),
	.D (n_4564),
	.CK (clk) );
   MX2X1 i_6180 ( .Y (n_4564),
	.S0 (n_5177),
	.B (pad_data_in[5]),
	.A (data_out[5]) );
   SDFFRHQX1 data_out_reg_6 ( .SI (data_out[5]),
	.SE (scan_en),
	.RN (n_4642),
	.Q (data_out[6]),
	.D (n_4570),
	.CK (clk) );
   MX2X1 i_6187 ( .Y (n_4570),
	.S0 (n_5177),
	.B (pad_data_in[6]),
	.A (data_out[6]) );
   NAND3BX1 i_26 ( .Y (n_28),
	.C (go),
	.B (bus_grant),
	.AN (read_cycle) );
   SDFFRHQX1 data_out_reg_7 ( .SI (data_out[6]),
	.SE (scan_en),
	.RN (n_4642),
	.Q (data_out[7]),
	.D (n_4576),
	.CK (clk) );
   MX2X1 i_6194 ( .Y (n_4576),
	.S0 (n_5177),
	.B (pad_data_in[7]),
	.A (data_out[7]) );
   SDFFRHQX1 data_out_reg_8 ( .SI (data_out[7]),
	.SE (FE_OFN135_scan_enI),
	.RN (n_4642),
	.Q (data_out[8]),
	.D (n_4582),
	.CK (clk) );
   MX2X1 i_6201 ( .Y (n_4582),
	.S0 (n_5177),
	.B (pad_data_in[8]),
	.A (data_out[8]) );
   SDFFRHQX1 data_out_reg_9 ( .SI (data_out[8]),
	.SE (FE_OFN19_scan_enI),
	.RN (n_4642),
	.Q (data_out[9]),
	.D (n_4588),
	.CK (clk) );
   MX2X1 i_6208 ( .Y (n_4588),
	.S0 (n_5177),
	.B (pad_data_in[9]),
	.A (data_out[9]) );
   AOI31X1 i_20 ( .Y (n_31),
	.B0 (present_state[1]),
	.A2 (go),
	.A1 (read_cycle),
	.A0 (bus_grant) );
   SDFFRHQX1 data_out_reg_10 ( .SI (data_out[9]),
	.SE (FE_OFN19_scan_enI),
	.RN (n_4642),
	.Q (data_out[10]),
	.D (n_4594),
	.CK (clk) );
   MX2X1 i_6215 ( .Y (n_4594),
	.S0 (n_5177),
	.B (pad_data_in[10]),
	.A (data_out[10]) );
   SDFFRHQX1 data_out_reg_11 ( .SI (data_out[10]),
	.SE (FE_OFN19_scan_enI),
	.RN (n_4642),
	.Q (data_out[11]),
	.D (n_4600),
	.CK (clk) );
   MX2X1 i_6222 ( .Y (n_4600),
	.S0 (n_5177),
	.B (pad_data_in[11]),
	.A (data_out[11]) );
   NOR3X1 i_0 ( .Y (n_5232),
	.C (n_4640),
	.B (present_state[1]),
	.A (present_state[0]) );
   SDFFRHQX1 data_out_reg_12 ( .SI (data_out[11]),
	.SE (FE_OFN19_scan_enI),
	.RN (n_4642),
	.Q (data_out[12]),
	.D (n_4606),
	.CK (clk) );
   MX2X1 i_6229 ( .Y (n_4606),
	.S0 (n_5177),
	.B (pad_data_in[12]),
	.A (data_out[12]) );
   NOR3BX1 i_19008 ( .Y (n_5226),
	.C (present_state[2]),
	.B (present_state[1]),
	.AN (present_state[0]) );
   SDFFRHQX1 data_out_reg_13 ( .SI (data_out[12]),
	.SE (FE_OFN19_scan_enI),
	.RN (n_4642),
	.Q (data_out[13]),
	.D (n_4612),
	.CK (clk) );
   MX2X1 i_6236 ( .Y (n_4612),
	.S0 (n_5177),
	.B (pad_data_in[13]),
	.A (data_out[13]) );
   AOI21X1 i_5 ( .Y (\nbus_626[0] ),
	.B0 (present_state[0]),
	.A1 (n_4640),
	.A0 (n_31) );
   SDFFRHQX1 data_out_reg_14 ( .SI (data_out[13]),
	.SE (FE_OFN19_scan_enI),
	.RN (n_4642),
	.Q (data_out[14]),
	.D (n_4618),
	.CK (clk) );
   MX2X1 i_6243 ( .Y (n_4618),
	.S0 (n_5177),
	.B (pad_data_in[14]),
	.A (data_out[14]) );
   AND2X1 i_7 ( .Y (n_5205),
	.B (present_state[1]),
	.A (present_state[0]) );
   SDFFRHQX1 data_out_reg_15 ( .SI (data_out[14]),
	.SE (FE_OFN19_scan_enI),
	.RN (n_4642),
	.Q (data_out[15]),
	.D (n_4624),
	.CK (clk) );
   MX2X1 i_6250 ( .Y (n_4624),
	.S0 (n_5177),
	.B (pad_data_in[15]),
	.A (data_out[15]) );
   NOR3BX1 i_9 ( .Y (n_5177),
	.C (present_state[2]),
	.B (present_state[0]),
	.AN (present_state[1]) );
   DFFRHQX1 write_reg ( .RN (n_4642),
	.Q (write),
	.D (n_5232),
	.CK (clk) );
   SDFFRHQX1 read_reg ( .SI (data_out[15]),
	.SE (FE_OFN6_scan_enI),
	.RN (n_4642),
	.Q (read),
	.D (n_5226),
	.CK (clk) );
   SDFFRHQX1 done_reg ( .SI (read),
	.SE (scan_en),
	.RN (n_4642),
	.Q (done),
	.D (n_5205),
	.CK (clk) );
   SDFFRHQX1 as_reg ( .SI (done),
	.SE (scan_en),
	.RN (n_4642),
	.Q (as),
	.D (n_21),
	.CK (clk) );
   SDFFRHQX1 bus_request_reg ( .SI (as),
	.SE (FE_OFN6_scan_enI),
	.RN (n_4642),
	.Q (bus_request),
	.D (n_21),
	.CK (clk) );
   INVX1 i_6322 ( .Y (n_4640),
	.A (present_state[2]) );
   INVX1 i_6323 ( .Y (n_4641),
	.A (n_23) );
   INVX1 i_6324 ( .Y (n_4642),
	.A (reset) );
   INVXL FE_OFC149_tdsp_data_out_15_ ( .Y (pad_data_out[15]),
	.A (FE_OFN149_tdsp_data_out_15_) );
   BUFX1 FE_OFC135_scan_enI ( .Y (FE_OFN135_scan_enI),
	.A (scan_en) );
   INVX2 FE_OFC111_t_addrs_0_ ( .Y (address[0]),
	.A (FE_OFN111_t_addrs_0_) );
   INVXL FE_OFC110_t_addrs_0_ ( .Y (FE_OFN111_t_addrs_0_),
	.A (FE_OFN110_t_addrs_0_) );
   INVX2 FE_OFC108_t_addrs_1_ ( .Y (address[1]),
	.A (FE_OFN108_t_addrs_1_) );
   INVXL FE_OFC107_t_addrs_1_ ( .Y (FE_OFN108_t_addrs_1_),
	.A (FE_OFN107_t_addrs_1_) );
   INVX2 FE_OFC105_t_addrs_2_ ( .Y (address[2]),
	.A (FE_OFN105_t_addrs_2_) );
   INVXL FE_OFC104_t_addrs_2_ ( .Y (FE_OFN105_t_addrs_2_),
	.A (FE_OFN104_t_addrs_2_) );
   INVX2 FE_OFC102_t_addrs_3_ ( .Y (address[3]),
	.A (FE_OFN102_t_addrs_3_) );
   INVXL FE_OFC101_t_addrs_3_ ( .Y (FE_OFN102_t_addrs_3_),
	.A (FE_OFN101_t_addrs_3_) );
   BUFX2 FE_OFC88_tdsp_data_out_0_ ( .Y (pad_data_out[0]),
	.A (FE_OFN88_tdsp_data_out_0_) );
   BUFX2 FE_OFC84_tdsp_data_out_1_ ( .Y (pad_data_out[1]),
	.A (FE_OFN84_tdsp_data_out_1_) );
   BUFX2 FE_OFC81_tdsp_data_out_2_ ( .Y (pad_data_out[2]),
	.A (FE_OFN81_tdsp_data_out_2_) );
   INVX2 FE_OFC77_tdsp_data_out_3_ ( .Y (pad_data_out[3]),
	.A (FE_OFN77_tdsp_data_out_3_) );
   INVXL FE_OFC76_tdsp_data_out_3_ ( .Y (FE_OFN77_tdsp_data_out_3_),
	.A (FE_OFN76_tdsp_data_out_3_) );
   INVX2 FE_OFC72_tdsp_data_out_4_ ( .Y (pad_data_out[4]),
	.A (FE_OFN72_tdsp_data_out_4_) );
   INVXL FE_OFC71_tdsp_data_out_4_ ( .Y (FE_OFN72_tdsp_data_out_4_),
	.A (FE_OFN71_tdsp_data_out_4_) );
   INVX2 FE_OFC67_tdsp_data_out_5_ ( .Y (pad_data_out[5]),
	.A (FE_OFN67_tdsp_data_out_5_) );
   INVXL FE_OFC66_tdsp_data_out_5_ ( .Y (FE_OFN67_tdsp_data_out_5_),
	.A (FE_OFN66_tdsp_data_out_5_) );
   INVX1 FE_OFC62_tdsp_data_out_6_ ( .Y (pad_data_out[6]),
	.A (FE_OFN62_tdsp_data_out_6_) );
   INVX1 FE_OFC57_tdsp_data_out_7_ ( .Y (pad_data_out[7]),
	.A (FE_OFN57_tdsp_data_out_7_) );
   INVX2 FE_OFC54_tdsp_data_out_8_ ( .Y (pad_data_out[8]),
	.A (FE_OFN54_tdsp_data_out_8_) );
   INVXL FE_OFC53_tdsp_data_out_8_ ( .Y (FE_OFN54_tdsp_data_out_8_),
	.A (FE_OFN53_tdsp_data_out_8_) );
   INVX2 FE_OFC48_tdsp_data_out_9_ ( .Y (pad_data_out[9]),
	.A (FE_OFN48_tdsp_data_out_9_) );
   INVXL FE_OFC44_tdsp_data_out_10_ ( .Y (pad_data_out[10]),
	.A (FE_OFN44_tdsp_data_out_10_) );
   INVXL FE_OFC40_tdsp_data_out_11_ ( .Y (pad_data_out[11]),
	.A (FE_OFN40_tdsp_data_out_11_) );
   INVX2 FE_OFC36_tdsp_data_out_12_ ( .Y (pad_data_out[12]),
	.A (FE_OFN36_tdsp_data_out_12_) );
   INVXL FE_OFC35_tdsp_data_out_12_ ( .Y (FE_OFN36_tdsp_data_out_12_),
	.A (FE_OFN35_tdsp_data_out_12_) );
   INVX2 FE_OFC31_tdsp_data_out_13_ ( .Y (pad_data_out[13]),
	.A (FE_OFN31_tdsp_data_out_13_) );
   INVXL FE_OFC30_tdsp_data_out_13_ ( .Y (FE_OFN31_tdsp_data_out_13_),
	.A (FE_OFN30_tdsp_data_out_13_) );
   INVXL FE_OFC25_tdsp_data_out_14_ ( .Y (pad_data_out[14]),
	.A (FE_OFN25_tdsp_data_out_14_) );
   BUFX16 FE_OFC22_tdsp_data_out_15_ ( .Y (FE_OFN149_tdsp_data_out_15_),
	.A (FE_OFN22_tdsp_data_out_15_) );
   BUFX1 FE_OFC19_scan_enI ( .Y (FE_OFN19_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC6_scan_enI ( .Y (FE_OFN6_scan_enI),
	.A (scan_en) );
endmodule

module decode_i (
	clk,
	reset,
	phi_1,
	phi_2,
	phi_3,
	phi_4,
	phi_5,
	phi_6,
	decode,
	p_data_out,
	ir,
	skip_one,
	read_prog,
	go_prog,
	read_data,
	go_data,
	read_port,
	go_port,
	decode_skip_one,
	scan_en,
	BG_scan_in,
	BG_scan_out );
   input clk;
   input reset;
   input phi_1;
   input phi_2;
   input phi_3;
   input phi_4;
   input phi_5;
   input phi_6;
   output [15:0] decode;
   input [15:0] p_data_out;
   output [15:0] ir;
   input skip_one;
   output read_prog;
   output go_prog;
   output read_data;
   output go_data;
   output read_port;
   output go_port;
   output decode_skip_one;
   input scan_en;
   input BG_scan_in;
   output BG_scan_out;

   // Internal wires
   wire \nbus_708[15] ;
   wire \nbus_669[15] ;
   wire n_73;
   wire n_140;
   wire n_4472;
   wire n_74;
   wire n_129;
   wire n_143;
   wire n_179;
   wire n_438;
   wire n_753;
   wire n_408;
   wire n_68;
   wire n_124;
   wire n_123;
   wire n_122;
   wire n_107;
   wire n_176;
   wire n_69;
   wire n_181;
   wire n_152;
   wire n_75;
   wire n_76;
   wire n_132;
   wire n_79;
   wire n_146;
   wire n_82;
   wire n_118;
   wire n_83;
   wire n_4473;
   wire n_84;
   wire n_150;
   wire n_161;
   wire n_135;
   wire n_88;
   wire n_145;
   wire n_90;
   wire n_139;
   wire n_163;
   wire n_165;
   wire n_134;
   wire n_92;
   wire n_564;
   wire n_141;
   wire n_4471;
   wire n_95;
   wire n_169;
   wire n_576;
   wire n_183;
   wire n_831;
   wire n_130;
   wire n_99;
   wire n_101;
   wire n_102;
   wire n_105;
   wire n_411;
   wire n_133;
   wire n_109;
   wire n_110;
   wire n_148;
   wire n_156;
   wire n_112;
   wire n_113;
   wire n_149;
   wire n_115;
   wire n_116;
   wire n_182;
   wire n_125;
   wire n_128;
   wire n_137;
   wire FE_OFN138_scan_enI;
   wire n_4225;
   wire n_4475;
   wire two_cycle;
   wire n_4228;
   wire n_4231;
   wire n_144;
   wire n_4237;
   wire n_4243;
   wire FE_OFN3_scan_enI;
   wire n_4249;
   wire n_4255;
   wire n_4261;
   wire n_4267;
   wire n_4273;
   wire n_151;
   wire FE_OFN134_scan_enI;
   wire n_4279;
   wire FE_OFN5_scan_enI;
   wire n_4285;
   wire n_4291;
   wire n_4297;
   wire n_155;
   wire n_4303;
   wire n_4309;
   wire n_4315;
   wire n_158;
   wire n_4321;
   wire FE_OFN168_scan_enI;
   wire n_4327;
   wire n_4333;
   wire n_4336;
   wire FE_OFN7_scan_enI;
   wire n_4339;
   wire n_4341;
   wire FE_OFN167_scan_enI;
   wire n_4345;
   wire n_4348;
   wire n_4351;
   wire n_4357;
   wire n_4363;
   wire FE_OFN169_scan_enI;
   wire n_4369;
   wire n_4375;
   wire n_4381;
   wire n_4387;
   wire n_4393;
   wire n_4399;
   wire n_4405;
   wire n_4411;
   wire n_174;
   wire n_4417;
   wire n_175;
   wire n_4423;
   wire FE_OFN170_scan_enI;
   wire n_4429;
   wire n_4435;
   wire n_4441;
   wire n_4447;
   wire n_4450;
   wire n_180;
   wire n_4453;
   wire n_4456;
   wire n_4474;
   wire n_4461;
   wire n_4459;
   wire n_4468;

   CLKBUFXL i_10028 ( .Y (ir[15]),
	.A (\nbus_708[15] ) );
   CLKBUFXL i_9919 ( .Y (decode[15]),
	.A (\nbus_669[15] ) );
   OAI21XL i_58 ( .Y (n_74),
	.B0 (n_4472),
	.A1 (n_140),
	.A0 (n_73) );
   NOR3X1 i_56 ( .Y (n_73),
	.C (n_143),
	.B (n_129),
	.A (decode[12]) );
   NOR2BX1 i_1036 ( .Y (n_438),
	.B (phi_3),
	.AN (n_179) );
   NOR2BX1 i_947 ( .Y (n_408),
	.B (phi_3),
	.AN (n_753) );
   AND2X1 i_574 ( .Y (n_753),
	.B (n_124),
	.A (n_68) );
   NAND4X1 i_35 ( .Y (n_69),
	.D (n_176),
	.C (n_107),
	.B (n_122),
	.A (n_123) );
   NAND2BX1 i_33 ( .Y (n_68),
	.B (decode_skip_one),
	.AN (n_181) );
   NAND2X1 i_61 ( .Y (n_75),
	.B (n_152),
	.A (decode[9]) );
   NAND3X1 i_62 ( .Y (n_76),
	.C (decode[11]),
	.B (decode[10]),
	.A (decode[8]) );
   NAND3X1 i_36 ( .Y (n_79),
	.C (n_75),
	.B (n_76),
	.A (n_132) );
   OAI21XL i_27 ( .Y (n_82),
	.B0 (decode[12]),
	.A1 (n_146),
	.A0 (decode[9]) );
   OAI21XL i_40 ( .Y (n_83),
	.B0 (n_118),
	.A1 (decode[11]),
	.A0 (decode[8]) );
   AOI211X1 i_74 ( .Y (n_84),
	.C0 (decode[15]),
	.B0 (decode[14]),
	.A1 (n_4473),
	.A0 (decode[13]) );
   NAND3X1 i_79 ( .Y (n_88),
	.C (n_135),
	.B (n_161),
	.A (n_150) );
   NOR4X1 i_82 ( .Y (n_90),
	.D (n_145),
	.C (decode[9]),
	.B (decode[11]),
	.A (decode[10]) );
   NAND4BBX1 i_34 ( .Y (n_92),
	.D (n_134),
	.C (n_165),
	.BN (n_163),
	.AN (n_139) );
   AOI21X1 i_1009 ( .Y (n_564),
	.B0 (phi_3),
	.A1 (n_4472),
	.A0 (n_92) );
   AOI22X1 i_25 ( .Y (n_95),
	.B1 (n_4471),
	.B0 (decode[11]),
	.A1 (n_141),
	.A0 (decode[10]) );
   OAI21XL i_808 ( .Y (n_576),
	.B0 (n_68),
	.A1 (n_169),
	.A0 (n_95) );
   OAI21XL i_570 ( .Y (n_831),
	.B0 (n_183),
	.A1 (n_124),
	.A0 (n_165) );
   NAND2X1 i_24 ( .Y (n_99),
	.B (n_130),
	.A (decode[11]) );
   OAI2BB1X1 i_31 ( .Y (n_101),
	.B0 (decode[13]),
	.A1N (n_99),
	.A0N (decode[14]) );
   NOR2X1 i_99 ( .Y (n_102),
	.B (decode[15]),
	.A (n_139) );
   AOI221X1 i_38 ( .Y (n_105),
	.C0 (n_102),
	.B1 (n_101),
	.B0 (decode[15]),
	.A1 (n_132),
	.A0 (decode[14]) );
   OAI21XL i_630 ( .Y (n_411),
	.B0 (n_68),
	.A1 (n_124),
	.A0 (n_105) );
   NAND3BX1 i_107 ( .Y (n_107),
	.C (n_143),
	.B (n_130),
	.AN (n_133) );
   NOR2X1 i_111 ( .Y (n_109),
	.B (n_4471),
	.A (decode[10]) );
   AOI21X1 i_112 ( .Y (n_110),
	.B0 (decode[11]),
	.A1 (n_141),
	.A0 (decode[10]) );
   NOR2BX1 i_113 ( .Y (n_112),
	.B (n_156),
	.AN (n_148) );
   AOI2BB1X1 i_114 ( .Y (n_113),
	.B0 (n_129),
	.A1N (n_109),
	.A0N (n_110) );
   AOI21X1 i_28 ( .Y (n_115),
	.B0 (decode[9]),
	.A1 (n_149),
	.A0 (n_146) );
   AOI31X1 i_30 ( .Y (n_116),
	.B0 (decode[13]),
	.A2 (decode[14]),
	.A1 (n_161),
	.A0 (n_150) );
   NAND2BX1 i_18 ( .Y (n_118),
	.B (decode[9]),
	.AN (n_149) );
   NAND2X1 i_118 ( .Y (n_122),
	.B (n_116),
	.A (decode[15]) );
   OAI21XL i_119 ( .Y (n_123),
	.B0 (decode[12]),
	.A1 (n_112),
	.A0 (n_113) );
   NAND2BX1 i_09006 ( .Y (n_124),
	.B (n_182),
	.AN (n_181) );
   NOR2BX1 i_23 ( .Y (n_125),
	.B (decode[14]),
	.AN (decode[13]) );
   NAND2X1 i_46 ( .Y (n_128),
	.B (decode[13]),
	.A (decode[14]) );
   NAND3X1 i_277 ( .Y (n_129),
	.C (decode[15]),
	.B (decode[13]),
	.A (decode[14]) );
   NOR2X1 i_346 ( .Y (n_130),
	.B (n_129),
	.A (decode[12]) );
   NAND3BX1 i_3 ( .Y (n_132),
	.C (decode[10]),
	.B (decode[8]),
	.AN (decode[9]) );
   NOR2BX1 i_17 ( .Y (n_133),
	.B (n_132),
	.AN (decode[11]) );
   AOI32X1 i_1 ( .Y (n_134),
	.B1 (n_133),
	.B0 (n_130),
	.A2 (decode[12]),
	.A1 (n_125),
	.A0 (decode[15]) );
   NOR2BX1 i_4 ( .Y (n_135),
	.B (decode[13]),
	.AN (decode[14]) );
   NOR4BX1 i_281 ( .Y (n_137),
	.D (decode[13]),
	.C (decode[12]),
	.B (decode[15]),
	.AN (decode[14]) );
   NOR3BX1 i_292 ( .Y (n_139),
	.C (decode[11]),
	.B (n_132),
	.AN (n_137) );
   NAND2BX1 i_12 ( .Y (n_140),
	.B (n_134),
	.AN (n_139) );
   NAND2X1 i_8 ( .Y (n_141),
	.B (decode[9]),
	.A (decode[8]) );
   SDFFRHQX1 two_cycle_reg ( .SI (BG_scan_in),
	.SE (FE_OFN138_scan_enI),
	.RN (n_4475),
	.Q (two_cycle),
	.D (n_4225),
	.CK (clk) );
   OAI211X1 i_5212 ( .Y (n_4225),
	.C0 (n_4228),
	.B0 (n_74),
	.A1 (n_438),
	.A0 (n_179) );
   NAND3X1 i_5214 ( .Y (n_4228),
	.C (two_cycle),
	.B (n_438),
	.A (n_74) );
   NAND4BXL i_48 ( .Y (n_143),
	.D (decode[9]),
	.C (decode[8]),
	.B (decode[10]),
	.AN (decode[11]) );
   SDFFRHQX1 decode_skip_one_reg ( .SI (two_cycle),
	.SE (scan_en),
	.RN (n_4475),
	.Q (decode_skip_one),
	.D (n_4231),
	.CK (clk) );
   MX2X1 i_5219 ( .Y (n_4231),
	.S0 (n_576),
	.B (n_182),
	.A (decode_skip_one) );
   NOR2BX1 i_67 ( .Y (n_144),
	.B (decode[15]),
	.AN (decode[12]) );
   SDFFRHQX1 decode_reg_0 ( .SI (decode_skip_one),
	.SE (scan_en),
	.RN (n_4475),
	.Q (decode[0]),
	.D (n_4237),
	.CK (clk) );
   MX2X1 i_5226 ( .Y (n_4237),
	.S0 (n_181),
	.B (decode[0]),
	.A (p_data_out[0]) );
   NAND2X1 i_422 ( .Y (n_145),
	.B (n_144),
	.A (n_125) );
   SDFFRHQX1 decode_reg_1 ( .SI (decode[0]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (decode[1]),
	.D (n_4243),
	.CK (clk) );
   MX2X1 i_5233 ( .Y (n_4243),
	.S0 (n_181),
	.B (decode[1]),
	.A (p_data_out[1]) );
   NAND2BX1 i_11 ( .Y (n_146),
	.B (decode[11]),
	.AN (decode[10]) );
   SDFFRHQX1 decode_reg_2 ( .SI (decode[1]),
	.SE (FE_OFN3_scan_enI),
	.RN (n_4475),
	.Q (decode[2]),
	.D (n_4249),
	.CK (clk) );
   MX2X1 i_5240 ( .Y (n_4249),
	.S0 (n_181),
	.B (decode[2]),
	.A (p_data_out[2]) );
   SDFFRHQX1 decode_reg_3 ( .SI (decode[2]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (decode[3]),
	.D (n_4255),
	.CK (clk) );
   MX2X1 i_5247 ( .Y (n_4255),
	.S0 (n_181),
	.B (decode[3]),
	.A (p_data_out[3]) );
   NOR2X1 i_269 ( .Y (n_148),
	.B (n_128),
	.A (decode[15]) );
   SDFFRHQX1 decode_reg_4 ( .SI (decode[3]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (decode[4]),
	.D (n_4261),
	.CK (clk) );
   MX2X1 i_5254 ( .Y (n_4261),
	.S0 (n_181),
	.B (decode[4]),
	.A (p_data_out[4]) );
   OR2X1 i_5 ( .Y (n_149),
	.B (decode[11]),
	.A (decode[10]) );
   SDFFRHQX1 decode_reg_5 ( .SI (decode[4]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (decode[5]),
	.D (n_4267),
	.CK (clk) );
   MX2X1 i_5261 ( .Y (n_4267),
	.S0 (n_181),
	.B (decode[5]),
	.A (p_data_out[5]) );
   NOR2X1 i_15 ( .Y (n_150),
	.B (n_149),
	.A (decode[12]) );
   SDFFRHQX1 decode_reg_6 ( .SI (decode[5]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (decode[6]),
	.D (n_4273),
	.CK (clk) );
   MX2X1 i_5268 ( .Y (n_4273),
	.S0 (n_181),
	.B (decode[6]),
	.A (p_data_out[6]) );
   NOR2BX1 i_22 ( .Y (n_151),
	.B (decode[12]),
	.AN (n_148) );
   SDFFSHQX1 decode_reg_7 ( .SN (n_4475),
	.SI (decode[6]),
	.SE (FE_OFN134_scan_enI),
	.Q (decode[7]),
	.D (n_4279),
	.CK (clk) );
   MX2X1 i_5275 ( .Y (n_4279),
	.S0 (n_181),
	.B (decode[7]),
	.A (p_data_out[7]) );
   NOR2X1 i_10 ( .Y (n_152),
	.B (decode[11]),
	.A (decode[8]) );
   SDFFSHQX1 decode_reg_8 ( .SN (n_4475),
	.SI (decode[7]),
	.SE (FE_OFN5_scan_enI),
	.Q (decode[8]),
	.D (n_4285),
	.CK (clk) );
   MX2X1 i_5282 ( .Y (n_4285),
	.S0 (n_181),
	.B (decode[8]),
	.A (p_data_out[8]) );
   SDFFSHQX1 decode_reg_9 ( .SN (n_4475),
	.SI (decode[8]),
	.SE (FE_OFN3_scan_enI),
	.Q (decode[9]),
	.D (n_4291),
	.CK (clk) );
   MX2X1 i_5289 ( .Y (n_4291),
	.S0 (n_181),
	.B (decode[9]),
	.A (p_data_out[9]) );
   SDFFSHQX1 decode_reg_10 ( .SN (n_4475),
	.SI (decode[9]),
	.SE (FE_OFN5_scan_enI),
	.Q (decode[10]),
	.D (n_4297),
	.CK (clk) );
   MX2X1 i_5296 ( .Y (n_4297),
	.S0 (n_181),
	.B (decode[10]),
	.A (p_data_out[10]) );
   AOI22X1 i_515 ( .Y (n_155),
	.B1 (n_150),
	.B0 (n_148),
	.A1 (n_79),
	.A0 (n_151) );
   SDFFSHQX1 decode_reg_11 ( .SN (n_4475),
	.SI (decode[10]),
	.SE (FE_OFN134_scan_enI),
	.Q (decode[11]),
	.D (n_4303),
	.CK (clk) );
   MX2X1 i_5303 ( .Y (n_4303),
	.S0 (n_181),
	.B (decode[11]),
	.A (p_data_out[11]) );
   AOI21X1 i_20 ( .Y (n_156),
	.B0 (n_146),
	.A1 (decode[9]),
	.A0 (decode[8]) );
   SDFFSHQX1 decode_reg_12 ( .SN (n_4475),
	.SI (decode[11]),
	.SE (scan_en),
	.Q (decode[12]),
	.D (n_4309),
	.CK (clk) );
   MX2X1 i_5310 ( .Y (n_4309),
	.S0 (n_181),
	.B (decode[12]),
	.A (p_data_out[12]) );
   SDFFSHQX1 decode_reg_13 ( .SN (n_4475),
	.SI (decode[12]),
	.SE (scan_en),
	.Q (decode[13]),
	.D (n_4315),
	.CK (clk) );
   MX2X1 i_5317 ( .Y (n_4315),
	.S0 (n_181),
	.B (decode[13]),
	.A (p_data_out[13]) );
   AOI32X1 i_77 ( .Y (n_158),
	.B1 (n_83),
	.B0 (n_137),
	.A2 (n_156),
	.A1 (n_148),
	.A0 (decode[12]) );
   SDFFSHQX1 decode_reg_14 ( .SN (n_4475),
	.SI (decode[13]),
	.SE (scan_en),
	.Q (decode[14]),
	.D (n_4321),
	.CK (clk) );
   MX2X1 i_5324 ( .Y (n_4321),
	.S0 (n_181),
	.B (decode[14]),
	.A (p_data_out[15]) );
   SDFFRHQX1 decode_reg_15 ( .SI (decode[14]),
	.SE (FE_OFN168_scan_enI),
	.RN (n_4475),
	.Q (\nbus_669[15] ),
	.D (n_4327),
	.CK (clk) );
   MX2X1 i_5331 ( .Y (n_4327),
	.S0 (n_181),
	.B (decode[15]),
	.A (p_data_out[14]) );
   SDFFRHQX1 go_port_reg ( .SI (\nbus_669[15] ),
	.SE (FE_OFN168_scan_enI),
	.RN (n_4475),
	.Q (go_port),
	.D (n_4333),
	.CK (clk) );
   OAI21XL i_5338 ( .Y (n_4333),
	.B0 (n_4336),
	.A1 (n_438),
	.A0 (n_179) );
   NAND2X1 i_5340 ( .Y (n_4336),
	.B (go_port),
	.A (n_438) );
   NOR2X1 i_9 ( .Y (n_161),
	.B (decode[9]),
	.A (decode[8]) );
   SDFFRHQX1 go_data_reg ( .SI (go_port),
	.SE (FE_OFN7_scan_enI),
	.RN (n_4475),
	.Q (go_data),
	.D (n_4339),
	.CK (clk) );
   OAI2BB1X1 i_5345 ( .Y (n_4339),
	.B0 (n_4341),
	.A1N (go_data),
	.A0N (n_564) );
   NAND2BX1 i_5346 ( .Y (n_4341),
	.B (n_831),
	.AN (n_564) );
   SDFFRHQX1 read_prog_reg ( .SI (go_data),
	.SE (FE_OFN167_scan_enI),
	.RN (n_4475),
	.Q (read_prog),
	.D (n_4345),
	.CK (clk) );
   OAI21XL i_5352 ( .Y (n_4345),
	.B0 (n_4348),
	.A1 (n_408),
	.A0 (n_753) );
   NAND2X1 i_5354 ( .Y (n_4348),
	.B (read_prog),
	.A (n_408) );
   NAND4BXL i_13 ( .Y (n_163),
	.D (n_88),
	.C (n_155),
	.B (n_158),
	.AN (n_84) );
   SDFFRHQX1 ir_reg_0 ( .SI (read_prog),
	.SE (scan_en),
	.RN (n_4475),
	.Q (ir[0]),
	.D (n_4351),
	.CK (clk) );
   MX2X1 i_5359 ( .Y (n_4351),
	.S0 (n_181),
	.B (ir[0]),
	.A (decode[0]) );
   SDFFRHQX1 ir_reg_1 ( .SI (ir[0]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (ir[1]),
	.D (n_4357),
	.CK (clk) );
   MX2X1 i_5366 ( .Y (n_4357),
	.S0 (n_181),
	.B (ir[1]),
	.A (decode[1]) );
   AOI21X1 i_14 ( .Y (n_165),
	.B0 (n_90),
	.A1 (n_144),
	.A0 (n_135) );
   SDFFRHQX1 ir_reg_2 ( .SI (ir[1]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (ir[2]),
	.D (n_4363),
	.CK (clk) );
   MX2X1 i_5373 ( .Y (n_4363),
	.S0 (n_181),
	.B (ir[2]),
	.A (decode[2]) );
   SDFFRHQX1 ir_reg_3 ( .SI (ir[2]),
	.SE (FE_OFN169_scan_enI),
	.RN (n_4475),
	.Q (ir[3]),
	.D (n_4369),
	.CK (clk) );
   MX2X1 i_5380 ( .Y (n_4369),
	.S0 (n_181),
	.B (ir[3]),
	.A (decode[3]) );
   SDFFRHQX1 ir_reg_4 ( .SI (ir[3]),
	.SE (FE_OFN169_scan_enI),
	.RN (n_4475),
	.Q (ir[4]),
	.D (n_4375),
	.CK (clk) );
   MX2X1 i_5387 ( .Y (n_4375),
	.S0 (n_181),
	.B (ir[4]),
	.A (decode[4]) );
   SDFFRHQX1 ir_reg_5 ( .SI (ir[4]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (ir[5]),
	.D (n_4381),
	.CK (clk) );
   MX2X1 i_5394 ( .Y (n_4381),
	.S0 (n_181),
	.B (ir[5]),
	.A (decode[5]) );
   NAND3BX1 i_92 ( .Y (n_169),
	.C (n_4472),
	.B (decode[12]),
	.AN (n_129) );
   SDFFRHQX1 ir_reg_6 ( .SI (ir[5]),
	.SE (scan_en),
	.RN (n_4475),
	.Q (ir[6]),
	.D (n_4387),
	.CK (clk) );
   MX2X1 i_5401 ( .Y (n_4387),
	.S0 (n_181),
	.B (ir[6]),
	.A (decode[6]) );
   SDFFSHQX1 ir_reg_7 ( .SN (n_4475),
	.SI (ir[6]),
	.SE (scan_en),
	.Q (ir[7]),
	.D (n_4393),
	.CK (clk) );
   MX2X1 i_5408 ( .Y (n_4393),
	.S0 (n_181),
	.B (ir[7]),
	.A (decode[7]) );
   SDFFSHQX2 ir_reg_8 ( .SN (n_4475),
	.SI (ir[7]),
	.SE (FE_OFN134_scan_enI),
	.Q (ir[8]),
	.D (n_4399),
	.CK (clk) );
   MX2X1 i_5415 ( .Y (n_4399),
	.S0 (n_181),
	.B (ir[8]),
	.A (decode[8]) );
   SDFFSHQX1 ir_reg_9 ( .SN (n_4475),
	.SI (ir[8]),
	.SE (scan_en),
	.Q (ir[9]),
	.D (n_4405),
	.CK (clk) );
   MX2X1 i_5422 ( .Y (n_4405),
	.S0 (n_181),
	.B (ir[9]),
	.A (decode[9]) );
   SDFFSHQX1 ir_reg_10 ( .SN (n_4475),
	.SI (ir[9]),
	.SE (scan_en),
	.Q (ir[10]),
	.D (n_4411),
	.CK (clk) );
   MX2X1 i_5429 ( .Y (n_4411),
	.S0 (n_181),
	.B (ir[10]),
	.A (decode[10]) );
   OAI211X1 i_122 ( .Y (n_174),
	.C0 (n_118),
	.B0 (n_137),
	.A1 (decode[11]),
	.A0 (decode[8]) );
   SDFFSHQX2 ir_reg_11 ( .SN (n_4475),
	.SI (ir[10]),
	.SE (scan_en),
	.Q (ir[11]),
	.D (n_4417),
	.CK (clk) );
   MX2X1 i_5436 ( .Y (n_4417),
	.S0 (n_181),
	.B (ir[11]),
	.A (decode[11]) );
   OAI22X1 i_123 ( .Y (n_175),
	.B1 (n_145),
	.B0 (n_115),
	.A1 (n_174),
	.A0 (n_139) );
   SDFFSHQX2 ir_reg_12 ( .SN (n_4475),
	.SI (ir[11]),
	.SE (FE_OFN168_scan_enI),
	.Q (ir[12]),
	.D (n_4423),
	.CK (clk) );
   MX2X1 i_5443 ( .Y (n_4423),
	.S0 (n_181),
	.B (ir[12]),
	.A (decode[12]) );
   AOI21X1 i_124 ( .Y (n_176),
	.B0 (n_175),
	.A1 (n_155),
	.A0 (n_151) );
   SDFFSHQX1 ir_reg_13 ( .SN (n_4475),
	.SI (ir[12]),
	.SE (FE_OFN170_scan_enI),
	.Q (ir[13]),
	.D (n_4429),
	.CK (clk) );
   MX2X1 i_5450 ( .Y (n_4429),
	.S0 (n_181),
	.B (ir[13]),
	.A (decode[13]) );
   SDFFSHQX1 ir_reg_14 ( .SN (n_4475),
	.SI (ir[13]),
	.SE (FE_OFN170_scan_enI),
	.Q (ir[14]),
	.D (n_4435),
	.CK (clk) );
   MX2X1 i_5457 ( .Y (n_4435),
	.S0 (n_181),
	.B (ir[14]),
	.A (decode[14]) );
   SDFFRHQX1 ir_reg_15 ( .SI (ir[14]),
	.SE (FE_OFN170_scan_enI),
	.RN (n_4475),
	.Q (\nbus_708[15] ),
	.D (n_4441),
	.CK (clk) );
   MX2X1 i_5464 ( .Y (n_4441),
	.S0 (n_181),
	.B (ir[15]),
	.A (decode[15]) );
   NAND4BXL i_401 ( .Y (n_179),
	.D (n_4472),
	.C (n_125),
	.B (decode[15]),
	.AN (decode[12]) );
   SDFFRHQX1 read_data_reg ( .SI (\nbus_708[15] ),
	.SE (FE_OFN7_scan_enI),
	.RN (n_4475),
	.Q (read_data),
	.D (n_4447),
	.CK (clk) );
   OAI21XL i_5471 ( .Y (n_4447),
	.B0 (n_4450),
	.A1 (n_564),
	.A0 (n_183) );
   NAND2X1 i_5473 ( .Y (n_4450),
	.B (read_data),
	.A (n_564) );
   NAND3BX1 i_663 ( .Y (n_180),
	.C (n_4475),
	.B (n_69),
	.AN (n_124) );
   SDFFRHQX1 read_port_reg ( .SI (read_data),
	.SE (FE_OFN7_scan_enI),
	.RN (n_4475),
	.Q (read_port),
	.D (n_4453),
	.CK (clk) );
   OAI21XL i_5478 ( .Y (n_4453),
	.B0 (n_4456),
	.A1 (n_438),
	.A0 (n_179) );
   NAND2X1 i_5480 ( .Y (n_4456),
	.B (read_port),
	.A (n_438) );
   NAND2BX1 i_2 ( .Y (n_181),
	.B (phi_6),
	.AN (skip_one) );
   SDFFRHQX1 go_prog_reg ( .SI (read_port),
	.SE (scan_en),
	.RN (n_4475),
	.Q (go_prog),
	.D (n_4474),
	.CK (clk) );
   AOI21X1 i_5485 ( .Y (n_4459),
	.B0 (n_4461),
	.A1 (go_prog),
	.A0 (n_408) );
   NOR2BX1 i_5486 ( .Y (n_4461),
	.B (n_408),
	.AN (n_411) );
   NOR2X1 i_21123 ( .Y (n_182),
	.B (two_cycle),
	.A (decode_skip_one) );
   SDFFHQX1 null_op_reg ( .SI (go_prog),
	.SE (FE_OFN167_scan_enI),
	.Q (BG_scan_out),
	.D (n_4468),
	.CK (clk) );
   AND2X1 i_5494 ( .Y (n_4468),
	.B (BG_scan_out),
	.A (n_180) );
   OAI21XL i_615 ( .Y (n_183),
	.B0 (n_4472),
	.A1 (n_163),
	.A0 (n_140) );
   INVX1 i_5659 ( .Y (n_4471),
	.A (n_161) );
   INVX1 i_5660 ( .Y (n_4472),
	.A (n_124) );
   INVX1 i_5661 ( .Y (n_4473),
	.A (n_82) );
   INVX1 i_5662 ( .Y (n_4474),
	.A (n_4459) );
   INVX1 i_5663 ( .Y (n_4475),
	.A (reset) );
   BUFX1 FE_OFC170_scan_enI ( .Y (FE_OFN170_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC169_scan_enI ( .Y (FE_OFN169_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC168_scan_enI ( .Y (FE_OFN168_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC167_scan_enI ( .Y (FE_OFN167_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC138_scan_enI ( .Y (FE_OFN138_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC134_scan_enI ( .Y (FE_OFN134_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC7_scan_enI ( .Y (FE_OFN7_scan_enI),
	.A (FE_OFN138_scan_enI) );
   BUFX1 FE_OFC5_scan_enI ( .Y (FE_OFN5_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC3_scan_enI ( .Y (FE_OFN3_scan_enI),
	.A (scan_en) );
endmodule

module execute_i (
	clk,
	reset,
	phi_1,
	phi_2,
	phi_3,
	phi_4,
	phi_5,
	phi_6,
	decode_skip_one,
	gez,
	gz,
	nz,
	z,
	lz,
	lez,
	ov,
	arnz,
	bioz,
	alu_result,
	mpy_result,
	mdr,
	pdr,
	ir,
	decode,
	ar,
	skip_one,
	fetch_branch,
	branch_stall,
	pc_acc,
	dmov_inc,
	dp,
	arp,
	ar0,
	ar1,
	pc,
	acc,
	p,
	top,
	alu_cmd,
	sel_op_a,
	sel_op_b,
	read_prog,
	go_prog,
	read_data,
	go_data,
	read_port,
	go_port,
	ovm,
	scan_en,
	BG_scan_in,
	BG_scan_out );
   input clk;
   input reset;
   input phi_1;
   input phi_2;
   input phi_3;
   input phi_4;
   input phi_5;
   input phi_6;
   input decode_skip_one;
   input gez;
   input gz;
   input nz;
   input z;
   input lz;
   input lez;
   output ov;
   input arnz;
   input bioz;
   input [32:0] alu_result;
   input [31:0] mpy_result;
   input [15:0] mdr;
   input [15:0] pdr;
   input [15:0] ir;
   input [15:0] decode;
   input [15:0] ar;
   output skip_one;
   output fetch_branch;
   output branch_stall;
   output pc_acc;
   output dmov_inc;
   output dp;
   output arp;
   output [15:0] ar0;
   output [15:0] ar1;
   output [15:0] pc;
   output [32:0] acc;
   output [31:0] p;
   output [15:0] top;
   output [3:0] alu_cmd;
   output [2:0] sel_op_a;
   output [2:0] sel_op_b;
   output read_prog;
   output go_prog;
   output read_data;
   output go_data;
   output read_port;
   output go_port;
   output ovm;
   input scan_en;
   input BG_scan_in;
   output BG_scan_out;

   // Internal wires
   wire [15:0] nbus_431;
   wire [2:0] nbus_435;
   wire [15:0] nbus_437;
   wire [2:0] nbus_439;
   wire n_7897;
   wire n_920;
   wire n_600;
   wire n_1031;
   wire n_595;
   wire n_718;
   wire n_1008;
   wire n_720;
   wire n_992;
   wire n_593;
   wire n_1006;
   wire n_590;
   wire n_794;
   wire n_850;
   wire n_792;
   wire n_855;
   wire n_4089;
   wire n_2082;
   wire n_585;
   wire n_474;
   wire \nbus_432[0] ;
   wire n_924;
   wire n_809;
   wire n_989;
   wire n_954;
   wire n_584;
   wire n_934;
   wire n_936;
   wire n_926;
   wire n_893;
   wire n_871;
   wire n_844;
   wire n_2534;
   wire n_828;
   wire n_4090;
   wire n_399;
   wire n_2610;
   wire n_896;
   wire n_580;
   wire n_578;
   wire n_576;
   wire n_573;
   wire n_571;
   wire n_966;
   wire n_570;
   wire n_568;
   wire n_566;
   wire n_967;
   wire n_565;
   wire n_563;
   wire n_561;
   wire n_968;
   wire n_560;
   wire n_558;
   wire n_556;
   wire n_969;
   wire n_555;
   wire n_553;
   wire n_551;
   wire n_970;
   wire n_550;
   wire n_548;
   wire n_546;
   wire n_971;
   wire n_545;
   wire n_543;
   wire n_541;
   wire n_972;
   wire n_540;
   wire n_538;
   wire n_536;
   wire n_973;
   wire n_535;
   wire n_533;
   wire n_531;
   wire n_974;
   wire n_529;
   wire n_528;
   wire n_526;
   wire n_975;
   wire n_524;
   wire n_523;
   wire n_982;
   wire n_519;
   wire n_518;
   wire n_516;
   wire n_984;
   wire n_513;
   wire n_511;
   wire n_981;
   wire n_508;
   wire n_506;
   wire n_978;
   wire three_cycle;
   wire n_2768;
   wire n_935;
   wire n_496;
   wire n_503;
   wire n_959;
   wire \nbus_428[0] ;
   wire \nbus_434[0] ;
   wire n_796;
   wire n_4082;
   wire n_952;
   wire n_811;
   wire n_960;
   wire n_497;
   wire n_499;
   wire n_380;
   wire n_879;
   wire n_940;
   wire n_922;
   wire n_829;
   wire n_804;
   wire n_955;
   wire n_950;
   wire n_494;
   wire n_820;
   wire n_951;
   wire n_948;
   wire n_949;
   wire n_941;
   wire n_491;
   wire n_2909;
   wire n_478;
   wire n_493;
   wire n_945;
   wire n_943;
   wire n_489;
   wire n_484;
   wire n_802;
   wire n_482;
   wire n_4080;
   wire n_788;
   wire n_481;
   wire n_485;
   wire n_912;
   wire n_913;
   wire n_483;
   wire n_889;
   wire n_863;
   wire n_800;
   wire n_475;
   wire \nbus_440[0] ;
   wire n_882;
   wire n_923;
   wire n_842;
   wire n_470;
   wire n_875;
   wire n_868;
   wire n_467;
   wire n_466;
   wire n_4220;
   wire n_464;
   wire n_910;
   wire n_3146;
   wire n_462;
   wire n_917;
   wire n_461;
   wire n_456;
   wire update_stall;
   wire n_1105;
   wire n_813;
   wire two_cycle;
   wire n_791;
   wire n_455;
   wire n_908;
   wire n_877;
   wire n_450;
   wire n_448;
   wire n_905;
   wire n_831;
   wire n_814;
   wire n_404;
   wire n_2765;
   wire n_446;
   wire n_4092;
   wire n_401;
   wire n_447;
   wire n_444;
   wire n_797;
   wire \nbus_436[0] ;
   wire n_839;
   wire n_440;
   wire n_836;
   wire n_442;
   wire n_835;
   wire n_438;
   wire n_899;
   wire n_4084;
   wire n_902;
   wire n_430;
   wire n_841;
   wire n_4085;
   wire n_432;
   wire n_843;
   wire n_431;
   wire n_429;
   wire branch_stall_delay;
   wire n_4083;
   wire n_2515;
   wire n_425;
   wire n_427;
   wire n_423;
   wire n_2384;
   wire n_805;
   wire n_890;
   wire n_823;
   wire n_886;
   wire n_883;
   wire n_424;
   wire n_1106;
   wire n_2115;
   wire n_414;
   wire n_830;
   wire n_2079;
   wire n_787;
   wire n_410;
   wire n_409;
   wire n_1940;
   wire n_784;
   wire n_395;
   wire n_790;
   wire n_851;
   wire n_383;
   wire n_407;
   wire n_406;
   wire n_405;
   wire n_403;
   wire n_2235;
   wire n_1833;
   wire n_816;
   wire n_793;
   wire n_400;
   wire n_396;
   wire n_697;
   wire n_1790;
   wire n_817;
   wire n_818;
   wire n_699;
   wire n_2387;
   wire n_4078;
   wire n_807;
   wire n_4077;
   wire n_795;
   wire n_1439;
   wire n_847;
   wire n_4079;
   wire n_382;
   wire n_869;
   wire n_722;
   wire n_724;
   wire n_1036;
   wire n_602;
   wire n_606;
   wire n_726;
   wire n_728;
   wire n_612;
   wire n_730;
   wire n_732;
   wire n_1018;
   wire n_614;
   wire n_619;
   wire n_734;
   wire n_736;
   wire n_1017;
   wire n_621;
   wire n_625;
   wire n_738;
   wire n_740;
   wire n_1033;
   wire n_627;
   wire n_631;
   wire n_742;
   wire n_744;
   wire n_4073;
   wire n_633;
   wire n_1015;
   wire n_635;
   wire n_637;
   wire n_748;
   wire n_747;
   wire n_1014;
   wire n_640;
   wire n_750;
   wire n_644;
   wire n_1044;
   wire n_1045;
   wire n_1013;
   wire n_647;
   wire n_754;
   wire n_651;
   wire n_1046;
   wire n_1047;
   wire n_4074;
   wire n_653;
   wire n_1012;
   wire n_655;
   wire n_758;
   wire n_658;
   wire n_1048;
   wire n_1049;
   wire n_1011;
   wire n_660;
   wire n_762;
   wire n_665;
   wire n_1050;
   wire n_1051;
   wire n_1010;
   wire n_668;
   wire n_766;
   wire n_672;
   wire n_1052;
   wire n_1053;
   wire n_1009;
   wire n_675;
   wire n_676;
   wire n_770;
   wire n_679;
   wire n_1054;
   wire n_1055;
   wire n_1056;
   wire n_1058;
   wire n_821;
   wire n_686;
   wire n_693;
   wire n_687;
   wire n_689;
   wire \nbus_430[0] ;
   wire n_1061;
   wire n_1943;
   wire n_1064;
   wire n_700;
   wire n_1793;
   wire n_925;
   wire n_937;
   wire n_1065;
   wire \nbus_429[2] ;
   wire n_932;
   wire \nbus_429[1] ;
   wire n_884;
   wire n_701;
   wire n_4100;
   wire n_872;
   wire n_704;
   wire n_806;
   wire n_705;
   wire n_962;
   wire \nbus_426[0] ;
   wire n_840;
   wire n_710;
   wire n_931;
   wire n_1076;
   wire n_712;
   wire n_4087;
   wire n_4086;
   wire n_713;
   wire n_808;
   wire n_714;
   wire n_715;
   wire n_716;
   wire n_717;
   wire n_1022;
   wire n_1086;
   wire n_1084;
   wire \nbus_425[15] ;
   wire n_1027;
   wire \nbus_425[14] ;
   wire n_4075;
   wire \nbus_425[13] ;
   wire n_1029;
   wire n_1025;
   wire n_1026;
   wire \nbus_425[12] ;
   wire n_1002;
   wire \nbus_425[11] ;
   wire n_4072;
   wire \nbus_425[10] ;
   wire n_1000;
   wire n_1001;
   wire \nbus_425[9] ;
   wire \nbus_425[8] ;
   wire n_999;
   wire n_751;
   wire \nbus_425[7] ;
   wire n_997;
   wire n_998;
   wire n_755;
   wire \nbus_425[6] ;
   wire n_759;
   wire \nbus_425[5] ;
   wire n_996;
   wire n_763;
   wire \nbus_425[4] ;
   wire n_994;
   wire n_995;
   wire n_767;
   wire \nbus_425[3] ;
   wire n_771;
   wire \nbus_425[2] ;
   wire n_1057;
   wire n_774;
   wire \nbus_425[1] ;
   wire n_837;
   wire n_777;
   wire n_780;
   wire n_782;
   wire \nbus_424[0] ;
   wire n_781;
   wire n_783;
   wire n_785;
   wire n_786;
   wire n_789;
   wire n_799;
   wire n_801;
   wire n_810;
   wire n_812;
   wire n_824;
   wire n_4088;
   wire n_832;
   wire n_838;
   wire update_it;
   wire n_856;
   wire n_859;
   wire n_864;
   wire n_865;
   wire n_873;
   wire n_876;
   wire n_880;
   wire n_895;
   wire n_897;
   wire n_914;
   wire n_915;
   wire n_4221;
   wire n_4076;
   wire n_927;
   wire n_928;
   wire n_930;
   wire n_4091;
   wire n_3104;
   wire n_1103;
   wire n_3107;
   wire FE_OFN163_scan_enI;
   wire n_3110;
   wire n_3113;
   wire n_3116;
   wire FE_OFN165_scan_enI;
   wire n_3122;
   wire FE_OFN9_scan_enI;
   wire n_4093;
   wire n_3130;
   wire n_3128;
   wire n_1114;
   wire n_1062;
   wire n_1111;
   wire n_3134;
   wire n_3137;
   wire n_3140;
   wire n_4094;
   wire n_3142;
   wire n_965;
   wire FE_OFN14_scan_enI;
   wire n_976;
   wire n_979;
   wire n_4101;
   wire n_3340;
   wire FE_OFN131_arp;
   wire n_1104;
   wire n_3343;
   wire FE_OFN139_scan_enI;
   wire n_3349;
   wire Q;
   wire n_3352;
   wire n_1108;
   wire n_4223;
   wire n_3354;
   wire n_3376;
   wire n_3379;
   wire n_3382;
   wire n_3385;
   wire n_3388;
   wire n_3394;
   wire n_3400;
   wire n_3406;
   wire FE_OFN166_scan_enI;
   wire n_3412;
   wire n_1005;
   wire n_3418;
   wire FE_OFN164_scan_enI;
   wire n_3424;
   wire n_3430;
   wire n_3436;
   wire n_3442;
   wire FE_OFN162_scan_enI;
   wire n_3448;
   wire n_3454;
   wire n_3460;
   wire n_3466;
   wire n_3472;
   wire n_3478;
   wire n_3484;
   wire n_3487;
   wire n_3490;
   wire n_1107;
   wire n_3493;
   wire n_1021;
   wire n_3514;
   wire n_3517;
   wire n_1028;
   wire FE_OFN142_scan_enI;
   wire n_1035;
   wire n_3616;
   wire FE_OFN129_dmov_inc;
   wire n_4081;
   wire n_3625;
   wire n_3631;
   wire n_3634;
   wire n_3637;
   wire n_1043;
   wire FE_OFN13_scan_enI;
   wire FE_OFN143_scan_enI;
   wire n_3736;
   wire n_3739;
   wire n_4095;
   wire n_3744;
   wire n_3742;
   wire n_4096;
   wire n_3750;
   wire n_3748;
   wire n_1071;
   wire n_3754;
   wire n_3757;
   wire n_4097;
   wire n_3769;
   wire FE_OFN17_scan_enI;
   wire n_1068;
   wire FE_OFN146_scan_enI;
   wire FE_OFN145_scan_enI;
   wire n_1081;
   wire FE_OFN171_scan_enI;
   wire n_3964;
   wire n_4222;
   wire n_3973;
   wire Q175;
   wire n_1109;
   wire n_4098;
   wire n_3978;
   wire n_3976;
   wire n_4099;
   wire n_1112;
   wire FE_OFN130_dmov_inc;

   INVXL i_10645 ( .Y (BG_scan_out),
	.A (n_7897) );
   INVXL i_10644 ( .Y (n_7897),
	.A (ar1[15]) );
   NAND2X1 i_579 ( .Y (n_600),
	.B (n_920),
	.A (mdr[14]) );
   NOR2X1 i_575 ( .Y (n_595),
	.B (n_1031),
	.A (ar[14]) );
   OAI221XL i_248240 ( .Y (nbus_431[15]),
	.C0 (n_593),
	.B1 (n_992),
	.B0 (n_720),
	.A1 (n_1008),
	.A0 (n_718) );
   NAND2X1 i_569 ( .Y (n_593),
	.B (n_920),
	.A (mdr[15]) );
   NOR2X1 i_567 ( .Y (n_590),
	.B (n_1006),
	.A (ar[15]) );
   AOI32X1 i_2507 ( .Y (n_2082),
	.B1 (n_4089),
	.B0 (n_855),
	.A2 (n_792),
	.A1 (n_850),
	.A0 (n_794) );
   NAND2X1 i_3501 ( .Y (\nbus_432[0] ),
	.B (n_474),
	.A (n_585) );
   NAND3BX1 i_551 ( .Y (n_585),
	.C (n_989),
	.B (n_809),
	.AN (n_924) );
   NAND2BX1 i_196 ( .Y (nbus_435[1]),
	.B (n_954),
	.AN (nbus_435[2]) );
   NAND4BXL i_195 ( .Y (nbus_435[2]),
	.D (n_926),
	.C (n_936),
	.B (n_934),
	.AN (n_584) );
   NOR3BX1 i_1694 ( .Y (n_584),
	.C (ir[14]),
	.B (ir[13]),
	.AN (ir[15]) );
   AOI32X1 i_2445 ( .Y (n_2534),
	.B1 (n_844),
	.B0 (mdr[0]),
	.A2 (n_871),
	.A1 (n_893),
	.A0 (ir[0]) );
   AOI31X1 i_2440 ( .Y (n_2610),
	.B0 (n_399),
	.A2 (n_4090),
	.A1 (n_828),
	.A0 (n_794) );
   OAI21XL i_398239 ( .Y (nbus_437[0]),
	.B0 (n_580),
	.A1 (pc[0]),
	.A0 (n_896) );
   NAND2X1 i_536 ( .Y (n_580),
	.B (n_896),
	.A (decode[0]) );
   OAI21XL i_388238 ( .Y (nbus_437[1]),
	.B0 (n_576),
	.A1 (n_578),
	.A0 (n_896) );
   XNOR2X1 i_244 ( .Y (n_578),
	.B (pc[0]),
	.A (pc[1]) );
   NAND2X1 i_532 ( .Y (n_576),
	.B (n_896),
	.A (decode[1]) );
   OAI21XL i_378237 ( .Y (nbus_437[2]),
	.B0 (n_571),
	.A1 (n_573),
	.A0 (n_896) );
   AOI21X1 i_243 ( .Y (n_573),
	.B0 (n_570),
	.A1 (n_966),
	.A0 (pc[2]) );
   NAND2X1 i_527 ( .Y (n_571),
	.B (n_896),
	.A (decode[2]) );
   NOR2X1 i_526 ( .Y (n_570),
	.B (n_966),
	.A (pc[2]) );
   OAI21XL i_368236 ( .Y (nbus_437[3]),
	.B0 (n_566),
	.A1 (n_568),
	.A0 (n_896) );
   AOI21X1 i_242 ( .Y (n_568),
	.B0 (n_565),
	.A1 (n_967),
	.A0 (pc[3]) );
   NAND2X1 i_522 ( .Y (n_566),
	.B (n_896),
	.A (decode[3]) );
   NOR2X1 i_521 ( .Y (n_565),
	.B (n_967),
	.A (pc[3]) );
   OAI21XL i_358235 ( .Y (nbus_437[4]),
	.B0 (n_561),
	.A1 (n_563),
	.A0 (n_896) );
   AOI21X1 i_241 ( .Y (n_563),
	.B0 (n_560),
	.A1 (n_968),
	.A0 (pc[4]) );
   NAND2X1 i_517 ( .Y (n_561),
	.B (n_896),
	.A (decode[4]) );
   NOR2X1 i_516 ( .Y (n_560),
	.B (n_968),
	.A (pc[4]) );
   OAI21XL i_348234 ( .Y (nbus_437[5]),
	.B0 (n_556),
	.A1 (n_558),
	.A0 (n_896) );
   AOI21X1 i_240 ( .Y (n_558),
	.B0 (n_555),
	.A1 (n_969),
	.A0 (pc[5]) );
   NAND2X1 i_512 ( .Y (n_556),
	.B (n_896),
	.A (decode[5]) );
   NOR2X1 i_511 ( .Y (n_555),
	.B (n_969),
	.A (pc[5]) );
   OAI21XL i_338233 ( .Y (nbus_437[6]),
	.B0 (n_551),
	.A1 (n_553),
	.A0 (n_896) );
   AOI21X1 i_239 ( .Y (n_553),
	.B0 (n_550),
	.A1 (n_970),
	.A0 (pc[6]) );
   NAND2X1 i_507 ( .Y (n_551),
	.B (n_896),
	.A (decode[6]) );
   NOR2X1 i_506 ( .Y (n_550),
	.B (n_970),
	.A (pc[6]) );
   OAI21XL i_32 ( .Y (nbus_437[7]),
	.B0 (n_546),
	.A1 (n_548),
	.A0 (n_896) );
   AOI21X1 i_238 ( .Y (n_548),
	.B0 (n_545),
	.A1 (n_971),
	.A0 (pc[7]) );
   NAND2X1 i_502 ( .Y (n_546),
	.B (n_896),
	.A (decode[7]) );
   NOR2X1 i_501 ( .Y (n_545),
	.B (n_971),
	.A (pc[7]) );
   OAI21XL i_318232 ( .Y (nbus_437[8]),
	.B0 (n_541),
	.A1 (n_543),
	.A0 (n_896) );
   AOI21X1 i_237 ( .Y (n_543),
	.B0 (n_540),
	.A1 (n_972),
	.A0 (pc[8]) );
   NAND2X1 i_497 ( .Y (n_541),
	.B (n_896),
	.A (decode[8]) );
   NOR2X1 i_496 ( .Y (n_540),
	.B (n_972),
	.A (pc[8]) );
   OAI21XL i_308231 ( .Y (nbus_437[9]),
	.B0 (n_536),
	.A1 (n_538),
	.A0 (n_896) );
   AOI21X1 i_236 ( .Y (n_538),
	.B0 (n_535),
	.A1 (n_973),
	.A0 (pc[9]) );
   NAND2X1 i_492 ( .Y (n_536),
	.B (n_896),
	.A (decode[9]) );
   NOR2X1 i_491 ( .Y (n_535),
	.B (n_973),
	.A (pc[9]) );
   OAI21XL i_298230 ( .Y (nbus_437[10]),
	.B0 (n_531),
	.A1 (n_533),
	.A0 (n_896) );
   AOI21X1 i_235 ( .Y (n_533),
	.B0 (n_529),
	.A1 (n_974),
	.A0 (pc[10]) );
   NAND2X1 i_487 ( .Y (n_531),
	.B (n_896),
	.A (decode[10]) );
   NOR2X1 i_485 ( .Y (n_529),
	.B (n_974),
	.A (pc[10]) );
   OAI21XL i_288229 ( .Y (nbus_437[11]),
	.B0 (n_526),
	.A1 (n_528),
	.A0 (n_896) );
   AOI21X1 i_234 ( .Y (n_528),
	.B0 (n_524),
	.A1 (n_975),
	.A0 (pc[11]) );
   NAND2X1 i_482 ( .Y (n_526),
	.B (n_896),
	.A (decode[11]) );
   NOR2X1 i_480 ( .Y (n_524),
	.B (n_975),
	.A (pc[11]) );
   MXI2X1 i_278228 ( .Y (nbus_437[12]),
	.S0 (n_896),
	.B (decode[12]),
	.A (n_523) );
   OAI31X1 i_233 ( .Y (n_523),
	.B0 (n_519),
	.A2 (pc[12]),
	.A1 (n_982),
	.A0 (n_973) );
   OAI21XL i_475 ( .Y (n_519),
	.B0 (pc[12]),
	.A1 (n_982),
	.A0 (n_973) );
   OAI21XL i_268227 ( .Y (nbus_437[13]),
	.B0 (n_516),
	.A1 (n_518),
	.A0 (n_896) );
   XNOR2X1 i_232 ( .Y (n_518),
	.B (n_984),
	.A (pc[13]) );
   NAND2X1 i_472 ( .Y (n_516),
	.B (n_896),
	.A (decode[13]) );
   OAI21XL i_258226 ( .Y (nbus_437[14]),
	.B0 (n_511),
	.A1 (n_513),
	.A0 (n_896) );
   XNOR2X1 i_231 ( .Y (n_513),
	.B (n_981),
	.A (pc[14]) );
   NAND2X1 i_467 ( .Y (n_511),
	.B (n_896),
	.A (decode[14]) );
   OAI21XL i_248225 ( .Y (nbus_437[15]),
	.B0 (n_506),
	.A1 (n_896),
	.A0 (n_508) );
   XNOR2X1 i_230 ( .Y (n_508),
	.B (n_978),
	.A (pc[15]) );
   NAND2X1 i_462 ( .Y (n_506),
	.B (n_896),
	.A (decode[15]) );
   NAND2X1 i_2796 ( .Y (n_2768),
	.B (three_cycle),
	.A (phi_6) );
   OR4X1 i_1818651 ( .Y (nbus_439[0]),
	.D (n_496),
	.C (n_935),
	.B (n_871),
	.A (n_584) );
   OAI21XL i_3732 ( .Y (\nbus_434[0] ),
	.B0 (\nbus_428[0] ),
	.A1 (n_959),
	.A0 (n_503) );
   AOI211X1 i_222 ( .Y (n_503),
	.C0 (n_584),
	.B0 (n_952),
	.A1 (n_4082),
	.A0 (n_796) );
   AOI211X1 i_185 ( .Y (\nbus_428[0] ),
	.C0 (n_499),
	.B0 (n_497),
	.A1 (n_960),
	.A0 (n_811) );
   AOI31X1 i_450 ( .Y (n_499),
	.B0 (n_959),
	.A2 (n_940),
	.A1 (n_879),
	.A0 (n_380) );
   NOR3X1 i_446 ( .Y (n_497),
	.C (n_804),
	.B (n_829),
	.A (n_922) );
   NAND4BXL i_1808650 ( .Y (nbus_439[1]),
	.D (n_954),
	.C (n_936),
	.B (n_950),
	.AN (n_955) );
   AND3X1 i_441 ( .Y (n_496),
	.C (n_829),
	.B (ir[14]),
	.A (ir[15]) );
   NAND2BX1 i_1798649 ( .Y (nbus_439[2]),
	.B (n_494),
	.AN (ir[15]) );
   OAI31X1 i_438 ( .Y (n_494),
	.B0 (ir[14]),
	.A2 (n_951),
	.A1 (n_820),
	.A0 (n_952) );
   AOI22X1 i_4078 ( .Y (n_2909),
	.B1 (n_491),
	.B0 (n_941),
	.A1 (n_949),
	.A0 (n_948) );
   AOI21X1 i_179 ( .Y (n_493),
	.B0 (n_478),
	.A1 (ir[4]),
	.A0 (ir[5]) );
   NAND4X1 i_221 ( .Y (n_491),
	.D (n_484),
	.C (n_489),
	.B (n_943),
	.A (n_945) );
   OAI21XL i_428 ( .Y (n_489),
	.B0 (n_4080),
	.A1 (n_482),
	.A0 (n_802) );
   OAI21XL i_178 ( .Y (n_485),
	.B0 (n_481),
	.A1 (n_788),
	.A0 (ir[9]) );
   NAND2X1 i_425 ( .Y (n_484),
	.B (n_912),
	.A (n_871) );
   AOI211X1 i_124 ( .Y (n_483),
	.C0 (n_913),
	.B0 (ir[10]),
	.A1 (ir[8]),
	.A0 (ir[9]) );
   NOR3X1 i_423 ( .Y (n_482),
	.C (n_483),
	.B (n_863),
	.A (n_889) );
   NAND2X1 i_422 ( .Y (n_481),
	.B (n_800),
	.A (ir[11]) );
   NOR2X1 i_419 ( .Y (n_478),
	.B (ir[4]),
	.A (ir[5]) );
   NAND2BX1 i_4136 ( .Y (\nbus_440[0] ),
	.B (n_474),
	.AN (n_475) );
   AOI21X1 i_416 ( .Y (n_475),
	.B0 (n_924),
	.A1 (n_882),
	.A0 (n_940) );
   NAND2X1 i_415 ( .Y (n_474),
	.B (n_811),
	.A (n_923) );
   NOR2X1 i_408 ( .Y (n_470),
	.B (n_842),
	.A (n_863) );
   NOR2BX1 i_404 ( .Y (n_467),
	.B (n_868),
	.AN (n_875) );
   AOI22X1 i_4206 ( .Y (n_3146),
	.B1 (n_910),
	.B0 (n_464),
	.A1 (n_4220),
	.A0 (n_466) );
   NAND2BX1 i_218 ( .Y (n_466),
	.B (n_462),
	.AN (n_920) );
   NAND4X1 i_219 ( .Y (n_464),
	.D (n_912),
	.C (n_456),
	.B (n_461),
	.A (n_917) );
   NAND3BX1 i_399 ( .Y (n_462),
	.C (n_1105),
	.B (phi_6),
	.AN (update_stall) );
   NAND2X1 i_389 ( .Y (n_461),
	.B (n_828),
	.A (three_cycle) );
   OAI21XL i_392 ( .Y (n_456),
	.B0 (n_809),
	.A1 (two_cycle),
	.A0 (n_813) );
   OAI221XL i_227 ( .Y (n_455),
	.C0 (n_800),
	.B1 (n_788),
	.B0 (n_791),
	.A1 (ir[10]),
	.A0 (ir[11]) );
   NAND3X1 i_380 ( .Y (n_450),
	.C (n_875),
	.B (n_877),
	.A (n_908) );
   OAI221XL i_3965 ( .Y (n_2765),
	.C0 (n_404),
	.B1 (n_814),
	.B0 (n_831),
	.A1 (n_905),
	.A0 (n_448) );
   AOI21X1 i_183 ( .Y (n_448),
	.B0 (n_828),
	.A1 (n_4092),
	.A0 (n_446) );
   OAI21XL i_79 ( .Y (n_447),
	.B0 (n_401),
	.A1 (n_829),
	.A0 (n_804) );
   NAND2X1 i_133 ( .Y (n_446),
	.B (n_804),
	.A (n_813) );
   OAI21XL i_3880 ( .Y (\nbus_436[0] ),
	.B0 (n_896),
	.A1 (n_797),
	.A0 (n_444) );
   AOI221X1 i_35 ( .Y (n_444),
	.C0 (n_442),
	.B1 (n_836),
	.B0 (n_440),
	.A1 (n_839),
	.A0 (ov) );
   NOR2BX1 i_367 ( .Y (n_442),
	.B (n_438),
	.AN (n_835) );
   OAI2BB1X1 i_248 ( .Y (n_440),
	.B0 (n_899),
	.A1N (n_791),
	.A0N (bioz) );
   AOI211X1 i_249 ( .Y (n_438),
	.C0 (n_430),
	.B0 (n_902),
	.A1 (n_4084),
	.A0 (gez) );
   NAND3X1 i_353 ( .Y (n_432),
	.C (lz),
	.B (n_4085),
	.A (n_841) );
   NAND3X1 i_354 ( .Y (n_431),
	.C (n_4085),
	.B (n_843),
	.A (lez) );
   NOR2BX1 i_351 ( .Y (n_430),
	.B (nz),
	.AN (n_844) );
   OR2X1 i_180 ( .Y (n_429),
	.B (n_844),
	.A (n_893) );
   AOI21X1 i_3737 ( .Y (n_2515),
	.B0 (n_4083),
	.A1 (branch_stall_delay),
	.A0 (phi_6) );
   AOI211X1 i_3576 ( .Y (n_2384),
	.C0 (n_423),
	.B0 (n_427),
	.A1 (n_425),
	.A0 (alu_result[32]) );
   AND4X1 i_343 ( .Y (n_427),
	.D (n_839),
	.C (ov),
	.B (n_794),
	.A (phi_1) );
   OAI2BB2X1 i_212 ( .Y (n_425),
	.B1 (n_890),
	.B0 (n_805),
	.A1N (n_4089),
	.A0N (n_811) );
   NAND4BXL i_213 ( .Y (n_424),
	.D (n_882),
	.C (n_883),
	.B (n_886),
	.AN (n_823) );
   AND4X1 i_341 ( .Y (n_423),
	.D (n_424),
	.C (alu_result[32]),
	.B (n_794),
	.A (phi_6) );
   NOR2X1 i_3659 ( .Y (n_2115),
	.B (phi_3),
	.A (n_1106) );
   AOI2BB1X1 i_3351 ( .Y (n_2079),
	.B0 (phi_3),
	.A1N (n_830),
	.A0N (n_414) );
   AOI21X1 i_210 ( .Y (n_414),
	.B0 (n_855),
	.A1 (n_792),
	.A0 (n_787) );
   NOR4BX1 i_3842 ( .Y (n_1940),
	.D (n_399),
	.C (phi_3),
	.B (n_409),
	.AN (n_410) );
   NAND2BX1 i_305 ( .Y (n_410),
	.B (n_395),
	.AN (n_784) );
   NOR2X1 i_302 ( .Y (n_409),
	.B (n_851),
	.A (n_790) );
   OAI211X1 i_295 ( .Y (n_407),
	.C0 (n_835),
	.B0 (n_794),
	.A1 (phi_1),
	.A0 (n_383) );
   NAND2X1 i_290 ( .Y (n_406),
	.B (n_835),
	.A (n_4085) );
   NOR4BX1 i_3157 ( .Y (n_1833),
	.D (n_2235),
	.C (n_403),
	.B (n_405),
	.AN (n_404) );
   NOR2X1 i_285 ( .Y (n_405),
	.B (n_830),
	.A (n_804) );
   NAND2X1 i_284 ( .Y (n_404),
	.B (n_447),
	.A (n_794) );
   AOI21X1 i_283 ( .Y (n_403),
	.B0 (n_830),
	.A1 (n_793),
	.A0 (n_816) );
   NAND2X1 i_280 ( .Y (n_401),
	.B (n_4090),
	.A (n_828) );
   OR2X1 i_3483 ( .Y (n_2235),
	.B (n_399),
	.A (n_400) );
   NOR2X1 i_275 ( .Y (n_400),
	.B (n_831),
	.A (n_814) );
   NOR2X1 i_274 ( .Y (n_399),
	.B (n_830),
	.A (n_813) );
   AOI222X1 i_3117 ( .Y (n_1790),
	.C1 (n_697),
	.C0 (n_796),
	.B1 (n_395),
	.B0 (n_396),
	.A1 (phi_1),
	.A0 (skip_one) );
   NAND3BX1 i_209 ( .Y (n_396),
	.C (n_699),
	.B (n_818),
	.AN (n_817) );
   AOI211X1 i_52 ( .Y (n_395),
	.C0 (branch_stall),
	.B0 (branch_stall_delay),
	.A1 (n_816),
	.A0 (n_793) );
   NAND2BX1 i_2462 ( .Y (nbus_435[0]),
	.B (n_2387),
	.AN (n_584) );
   AOI211X1 i_2797 ( .Y (n_2387),
	.C0 (n_802),
	.B0 (n_807),
	.A1 (n_4078),
	.A0 (ir[14]) );
   OAI32X1 i_2874 ( .Y (n_1439),
	.B1 (n_795),
	.B0 (n_784),
	.A2 (n_4077),
	.A1 (n_793),
	.A0 (n_797) );
   NOR3BX1 i_1731 ( .Y (n_383),
	.C (n_836),
	.B (n_839),
	.AN (n_847) );
   NAND2BX1 i_63 ( .Y (n_382),
	.B (n_4079),
	.AN (n_913) );
   NAND3X1 i_2232 ( .Y (n_380),
	.C (n_869),
	.B (ir[0]),
	.A (ir[2]) );
   OAI221XL i_258241 ( .Y (nbus_431[14]),
	.C0 (n_600),
	.B1 (n_992),
	.B0 (n_724),
	.A1 (n_1008),
	.A0 (n_722) );
   NOR2X1 i_586 ( .Y (n_602),
	.B (n_1036),
	.A (ar[13]) );
   NAND2X1 i_589 ( .Y (n_606),
	.B (n_920),
	.A (mdr[13]) );
   OAI221XL i_268242 ( .Y (nbus_431[13]),
	.C0 (n_606),
	.B1 (n_992),
	.B0 (n_728),
	.A1 (n_1008),
	.A0 (n_726) );
   NAND2X1 i_597 ( .Y (n_612),
	.B (n_920),
	.A (mdr[12]) );
   OAI221XL i_278243 ( .Y (nbus_431[12]),
	.C0 (n_612),
	.B1 (n_992),
	.B0 (n_732),
	.A1 (n_1008),
	.A0 (n_730) );
   NOR2X1 i_602 ( .Y (n_614),
	.B (n_1018),
	.A (ar[11]) );
   NAND2X1 i_606 ( .Y (n_619),
	.B (n_920),
	.A (mdr[11]) );
   OAI221XL i_288244 ( .Y (nbus_431[11]),
	.C0 (n_619),
	.B1 (n_992),
	.B0 (n_736),
	.A1 (n_1008),
	.A0 (n_734) );
   NOR2X1 i_611 ( .Y (n_621),
	.B (n_1017),
	.A (ar[10]) );
   NAND2X1 i_614 ( .Y (n_625),
	.B (n_920),
	.A (mdr[10]) );
   OAI221XL i_298245 ( .Y (nbus_431[10]),
	.C0 (n_625),
	.B1 (n_992),
	.B0 (n_740),
	.A1 (n_1008),
	.A0 (n_738) );
   NOR2X1 i_619 ( .Y (n_627),
	.B (n_1033),
	.A (ar[9]) );
   NAND2X1 i_622 ( .Y (n_631),
	.B (n_920),
	.A (mdr[9]) );
   OAI221XL i_308246 ( .Y (nbus_431[9]),
	.C0 (n_631),
	.B1 (n_992),
	.B0 (n_744),
	.A1 (n_1008),
	.A0 (n_742) );
   OAI21XL i_627 ( .Y (n_633),
	.B0 (ar[8]),
	.A1 (ar[7]),
	.A0 (n_4073) );
   NOR2X1 i_629 ( .Y (n_635),
	.B (n_1015),
	.A (ar[8]) );
   NAND2X1 i_630 ( .Y (n_637),
	.B (n_920),
	.A (mdr[8]) );
   OAI221XL i_318247 ( .Y (nbus_431[8]),
	.C0 (n_637),
	.B1 (n_992),
	.B0 (n_747),
	.A1 (n_1008),
	.A0 (n_748) );
   NOR2X1 i_636 ( .Y (n_640),
	.B (n_1014),
	.A (ar[7]) );
   NOR2X1 i_640 ( .Y (n_644),
	.B (n_1008),
	.A (n_750) );
   NAND2X1 i_328248 ( .Y (nbus_431[7]),
	.B (n_1045),
	.A (n_1044) );
   NOR2X1 i_645 ( .Y (n_647),
	.B (n_1013),
	.A (ar[6]) );
   NOR2X1 i_649 ( .Y (n_651),
	.B (n_1008),
	.A (n_754) );
   NAND2X1 i_338249 ( .Y (nbus_431[6]),
	.B (n_1047),
	.A (n_1046) );
   OAI21XL i_653 ( .Y (n_653),
	.B0 (ar[5]),
	.A1 (ar[4]),
	.A0 (n_4074) );
   NOR2X1 i_655 ( .Y (n_655),
	.B (n_1012),
	.A (ar[5]) );
   NOR2X1 i_658 ( .Y (n_658),
	.B (n_992),
	.A (n_758) );
   NAND2X1 i_348250 ( .Y (nbus_431[5]),
	.B (n_1049),
	.A (n_1048) );
   NOR2X1 i_662 ( .Y (n_660),
	.B (n_1011),
	.A (ar[4]) );
   NOR2X1 i_667 ( .Y (n_665),
	.B (n_1008),
	.A (n_762) );
   NAND2X1 i_358251 ( .Y (nbus_431[4]),
	.B (n_1051),
	.A (n_1050) );
   NOR2X1 i_672 ( .Y (n_668),
	.B (n_1010),
	.A (ar[3]) );
   NOR2X1 i_676 ( .Y (n_672),
	.B (n_1008),
	.A (n_766) );
   NAND2X1 i_368252 ( .Y (nbus_431[3]),
	.B (n_1053),
	.A (n_1052) );
   NOR2X1 i_681 ( .Y (n_675),
	.B (ar[2]),
	.A (n_1009) );
   OAI21XL i_682 ( .Y (n_676),
	.B0 (ar[2]),
	.A1 (ar[1]),
	.A0 (ar[0]) );
   NOR2X1 i_685 ( .Y (n_679),
	.B (n_1008),
	.A (n_770) );
   NAND2X1 i_378253 ( .Y (nbus_431[2]),
	.B (n_1055),
	.A (n_1054) );
   NAND2X1 i_388254 ( .Y (nbus_431[1]),
	.B (n_1058),
	.A (n_1056) );
   NAND4X1 i_696 ( .Y (n_686),
	.D (n_4079),
	.C (n_821),
	.B (ir[12]),
	.A (ir[11]) );
   NAND2BX1 i_699 ( .Y (n_687),
	.B (n_948),
	.AN (n_693) );
   OAI21XL i_223 ( .Y (n_689),
	.B0 (n_686),
	.A1 (n_4080),
	.A0 (n_863) );
   OAI2BB1X1 i_3282 ( .Y (\nbus_430[0] ),
	.B0 (n_687),
	.A1N (n_941),
	.A0N (n_689) );
   AND2X1 i_136 ( .Y (n_693),
	.B (n_992),
	.A (n_1008) );
   OAI21XL i_398255 ( .Y (nbus_431[0]),
	.B0 (n_1061),
	.A1 (ar[0]),
	.A0 (n_693) );
   NOR2BX1 i_2655 ( .Y (n_1943),
	.B (n_409),
	.AN (n_2610) );
   OAI22X1 i_76 ( .Y (n_697),
	.B1 (n_805),
	.B0 (n_804),
	.A1 (n_4220),
	.A0 (n_814) );
   NAND2X1 i_55 ( .Y (n_699),
	.B (three_cycle),
	.A (phi_4) );
   AOI22X1 i_228 ( .Y (n_700),
	.B1 (n_830),
	.B0 (n_1064),
	.A1 (n_793),
	.A0 (n_816) );
   AOI22X1 i_2385 ( .Y (n_1793),
	.B1 (n_796),
	.B0 (n_697),
	.A1 (n_699),
	.A0 (n_700) );
   OR3XL i_1798667 ( .Y (\nbus_429[2] ),
	.C (n_1065),
	.B (n_937),
	.A (n_925) );
   NOR4BX1 i_1808668 ( .Y (\nbus_429[1] ),
	.D (n_932),
	.C (n_937),
	.B (n_821),
	.AN (n_926) );
   NAND2X1 i_722 ( .Y (n_701),
	.B (n_884),
	.A (n_809) );
   NOR3X1 i_203 ( .Y (n_704),
	.C (n_872),
	.B (n_4100),
	.A (ir[10]) );
   AOI21X1 i_726 ( .Y (n_705),
	.B0 (n_806),
	.A1 (n_701),
	.A0 (n_872) );
   OAI32X1 i_2924 ( .Y (\nbus_426[0] ),
	.B1 (n_962),
	.B0 (n_924),
	.A2 (n_804),
	.A1 (n_818),
	.A0 (n_922) );
   AOI21X1 i_73 ( .Y (n_710),
	.B0 (n_840),
	.A1 (n_806),
	.A0 (n_788) );
   NOR2X1 i_747 ( .Y (n_712),
	.B (n_1076),
	.A (n_931) );
   OAI32X1 i_112 ( .Y (n_713),
	.B1 (n_4086),
	.B0 (n_710),
	.A2 (n_4087),
	.A1 (n_844),
	.A0 (n_841) );
   OAI21XL i_743 ( .Y (n_714),
	.B0 (ir[12]),
	.A1 (n_808),
	.A0 (n_821) );
   NAND2X1 i_744 ( .Y (n_715),
	.B (n_4080),
	.A (n_802) );
   NAND3BX1 i_745 ( .Y (n_716),
	.C (n_813),
	.B (n_809),
	.AN (n_989) );
   NOR3X1 i_746 ( .Y (n_717),
	.C (n_863),
	.B (n_951),
	.A (n_935) );
   XNOR2X1 i_83 ( .Y (n_718),
	.B (n_1022),
	.A (ar[15]) );
   AOI21X1 i_84 ( .Y (n_720),
	.B0 (n_590),
	.A1 (n_1006),
	.A0 (ar[15]) );
   OAI221XL i_248256 ( .Y (\nbus_425[15] ),
	.C0 (n_593),
	.B1 (n_720),
	.B0 (n_1084),
	.A1 (n_718),
	.A0 (n_1086) );
   AOI21X1 i_85 ( .Y (n_722),
	.B0 (n_595),
	.A1 (n_1031),
	.A0 (ar[14]) );
   XNOR2X1 i_86 ( .Y (n_724),
	.B (n_1027),
	.A (ar[14]) );
   OAI221XL i_258257 ( .Y (\nbus_425[14] ),
	.C0 (n_600),
	.B1 (n_724),
	.B0 (n_1084),
	.A1 (n_722),
	.A0 (n_1086) );
   AOI21X1 i_87 ( .Y (n_726),
	.B0 (n_602),
	.A1 (n_1036),
	.A0 (ar[13]) );
   AOI21X1 i_88 ( .Y (n_728),
	.B0 (n_1027),
	.A1 (n_4075),
	.A0 (ar[13]) );
   OAI221XL i_268258 ( .Y (\nbus_425[13] ),
	.C0 (n_606),
	.B1 (n_1084),
	.B0 (n_728),
	.A1 (n_726),
	.A0 (n_1086) );
   XNOR2X1 i_89 ( .Y (n_730),
	.B (n_1029),
	.A (ar[12]) );
   AOI21X1 i_90 ( .Y (n_732),
	.B0 (n_1026),
	.A1 (n_1025),
	.A0 (ar[12]) );
   OAI221XL i_278259 ( .Y (\nbus_425[12] ),
	.C0 (n_612),
	.B1 (n_732),
	.B0 (n_1084),
	.A1 (n_730),
	.A0 (n_1086) );
   AOI21X1 i_91 ( .Y (n_734),
	.B0 (n_614),
	.A1 (n_1018),
	.A0 (ar[11]) );
   XNOR2X1 i_92 ( .Y (n_736),
	.B (n_1002),
	.A (ar[11]) );
   OAI221XL i_288260 ( .Y (\nbus_425[11] ),
	.C0 (n_619),
	.B1 (n_736),
	.B0 (n_1084),
	.A1 (n_734),
	.A0 (n_1086) );
   AOI21X1 i_93 ( .Y (n_738),
	.B0 (n_621),
	.A1 (n_1017),
	.A0 (ar[10]) );
   AOI21X1 i_94 ( .Y (n_740),
	.B0 (n_1002),
	.A1 (n_4072),
	.A0 (ar[10]) );
   OAI221XL i_298261 ( .Y (\nbus_425[10] ),
	.C0 (n_625),
	.B1 (n_1084),
	.B0 (n_740),
	.A1 (n_738),
	.A0 (n_1086) );
   AOI21X1 i_95 ( .Y (n_742),
	.B0 (n_627),
	.A1 (n_1033),
	.A0 (ar[9]) );
   AOI21X1 i_96 ( .Y (n_744),
	.B0 (n_1001),
	.A1 (n_1000),
	.A0 (ar[9]) );
   OAI221XL i_308262 ( .Y (\nbus_425[9] ),
	.C0 (n_631),
	.B1 (n_744),
	.B0 (n_1084),
	.A1 (n_742),
	.A0 (n_1086) );
   AND2X1 i_97 ( .Y (n_747),
	.B (n_633),
	.A (n_1000) );
   AOI21X1 i_106 ( .Y (n_748),
	.B0 (n_635),
	.A1 (n_1015),
	.A0 (ar[8]) );
   OAI221XL i_318263 ( .Y (\nbus_425[8] ),
	.C0 (n_637),
	.B1 (n_1084),
	.B0 (n_747),
	.A1 (n_748),
	.A0 (n_1086) );
   AOI21X1 i_99 ( .Y (n_750),
	.B0 (n_640),
	.A1 (n_1014),
	.A0 (ar[7]) );
   AOI21X1 i_100 ( .Y (n_751),
	.B0 (n_999),
	.A1 (n_4073),
	.A0 (ar[7]) );
   OAI221XL i_328264 ( .Y (\nbus_425[7] ),
	.C0 (n_1044),
	.B1 (n_750),
	.B0 (n_1086),
	.A1 (n_1084),
	.A0 (n_751) );
   AOI21X1 i_101 ( .Y (n_754),
	.B0 (n_647),
	.A1 (n_1013),
	.A0 (ar[6]) );
   AOI21X1 i_120 ( .Y (n_755),
	.B0 (n_998),
	.A1 (n_997),
	.A0 (ar[6]) );
   OAI221XL i_338265 ( .Y (\nbus_425[6] ),
	.C0 (n_1046),
	.B1 (n_754),
	.B0 (n_1086),
	.A1 (n_755),
	.A0 (n_1084) );
   AND2X1 i_102 ( .Y (n_758),
	.B (n_653),
	.A (n_997) );
   AOI21X1 i_109 ( .Y (n_759),
	.B0 (n_655),
	.A1 (n_1012),
	.A0 (ar[5]) );
   OAI221XL i_348266 ( .Y (\nbus_425[5] ),
	.C0 (n_1048),
	.B1 (n_1084),
	.B0 (n_758),
	.A1 (n_759),
	.A0 (n_1086) );
   AOI21X1 i_103 ( .Y (n_762),
	.B0 (n_660),
	.A1 (n_1011),
	.A0 (ar[4]) );
   AOI21X1 i_121 ( .Y (n_763),
	.B0 (n_996),
	.A1 (n_4074),
	.A0 (ar[4]) );
   OAI221XL i_358267 ( .Y (\nbus_425[4] ),
	.C0 (n_1050),
	.B1 (n_762),
	.B0 (n_1086),
	.A1 (n_1084),
	.A0 (n_763) );
   AOI21X1 i_110 ( .Y (n_766),
	.B0 (n_668),
	.A1 (n_1010),
	.A0 (ar[3]) );
   AOI21X1 i_125 ( .Y (n_767),
	.B0 (n_995),
	.A1 (n_994),
	.A0 (ar[3]) );
   OAI221XL i_368268 ( .Y (\nbus_425[3] ),
	.C0 (n_1052),
	.B1 (n_766),
	.B0 (n_1086),
	.A1 (n_767),
	.A0 (n_1084) );
   AOI21X1 i_104 ( .Y (n_770),
	.B0 (n_675),
	.A1 (n_1009),
	.A0 (ar[2]) );
   AND2X1 i_122 ( .Y (n_771),
	.B (n_676),
	.A (n_994) );
   OAI221XL i_378269 ( .Y (\nbus_425[2] ),
	.C0 (n_1054),
	.B1 (n_770),
	.B0 (n_1086),
	.A1 (n_1084),
	.A0 (n_771) );
   NAND2BX1 i_824 ( .Y (n_774),
	.B (n_1057),
	.AN (n_1084) );
   OAI211X1 i_388270 ( .Y (\nbus_425[1] ),
	.C0 (n_774),
	.B0 (n_1056),
	.A1 (n_1057),
	.A0 (n_1086) );
   NAND4BXL i_829 ( .Y (n_777),
	.D (n_821),
	.C (ir[12]),
	.B (ir[11]),
	.AN (n_837) );
   OAI31X1 i_225 ( .Y (n_780),
	.B0 (n_777),
	.A2 (n_863),
	.A1 (n_837),
	.A0 (ir[11]) );
   AOI22X1 i_2811 ( .Y (\nbus_424[0] ),
	.B1 (n_948),
	.B0 (n_782),
	.A1 (n_941),
	.A0 (n_780) );
   NAND2BX1 i_834 ( .Y (n_781),
	.B (n_782),
	.AN (ar[0]) );
   NAND2X1 i_137 ( .Y (n_782),
	.B (n_1084),
	.A (n_1086) );
   NOR2X1 i_71 ( .Y (n_783),
	.B (n_4092),
	.A (three_cycle) );
   NAND2X1 i_21022 ( .Y (n_784),
	.B (n_783),
	.A (phi_6) );
   NAND2X1 i_38 ( .Y (n_785),
	.B (ir[14]),
	.A (ir[15]) );
   NAND3X1 i_78 ( .Y (n_786),
	.C (ir[13]),
	.B (ir[14]),
	.A (ir[15]) );
   NOR2X1 i_1701 ( .Y (n_787),
	.B (n_786),
	.A (ir[12]) );
   NAND2X1 i_23 ( .Y (n_788),
	.B (ir[8]),
	.A (ir[10]) );
   NOR2X1 i_28 ( .Y (n_789),
	.B (n_788),
	.A (ir[9]) );
   NAND2X1 i_115 ( .Y (n_790),
	.B (n_789),
	.A (ir[11]) );
   NOR2BX1 i_20 ( .Y (n_791),
	.B (ir[11]),
	.AN (ir[9]) );
   NOR2BX1 i_193 ( .Y (n_792),
	.B (n_788),
	.AN (n_791) );
   OAI21XL i_0 ( .Y (n_793),
	.B0 (n_787),
	.A1 (n_4084),
	.A0 (n_792) );
   NOR2X1 i_29 ( .Y (n_794),
	.B (branch_stall),
	.A (branch_stall_delay) );
   NAND2BX1 i_189 ( .Y (n_795),
	.B (n_794),
	.AN (n_793) );
   NOR2X1 i_44 ( .Y (n_796),
	.B (two_cycle),
	.A (three_cycle) );
   NAND2X1 i_170 ( .Y (n_797),
	.B (phi_1),
	.A (n_794) );
   NOR2X1 i_62 ( .Y (n_799),
	.B (ir[9]),
	.A (ir[10]) );
   NAND2X1 i_21 ( .Y (n_800),
	.B (n_4100),
	.A (n_799) );
   NOR2X1 i_37 ( .Y (n_801),
	.B (n_800),
	.A (ir[11]) );
   NOR2X1 i_1765 ( .Y (n_802),
	.B (n_785),
	.A (ir[13]) );
   NAND3BX1 i_22 ( .Y (n_804),
	.C (n_801),
	.B (n_802),
	.AN (ir[12]) );
   NAND2X1 i_67 ( .Y (n_805),
	.B (n_794),
	.A (phi_3) );
   NAND2X1 i_24 ( .Y (n_806),
	.B (n_4100),
	.A (ir[10]) );
   NOR2X1 i_256 ( .Y (n_807),
	.B (ir[13]),
	.A (ir[15]) );
   AND2X1 i_1756 ( .Y (n_808),
	.B (n_807),
	.A (ir[14]) );
   NOR2BX1 i_1790 ( .Y (n_809),
	.B (ir[12]),
	.AN (n_808) );
   AND2X1 i_194 ( .Y (n_810),
	.B (n_791),
	.A (n_809) );
   AND2X1 i_1845 ( .Y (n_811),
	.B (n_4087),
	.A (n_810) );
   NOR3X1 i_45 ( .Y (n_812),
	.C (ir[11]),
	.B (n_788),
	.A (ir[9]) );
   AOI21X1 i_1808 ( .Y (n_813),
	.B0 (n_811),
	.A1 (n_812),
	.A0 (n_809) );
   NAND2BX1 i_200 ( .Y (n_814),
	.B (n_794),
	.AN (n_813) );
   NAND3BX1 i_1763 ( .Y (n_816),
	.C (ir[13]),
	.B (ir[15]),
	.AN (ir[14]) );
   AOI21X1 i_27 ( .Y (n_817),
	.B0 (n_4220),
	.A1 (three_cycle),
	.A0 (two_cycle) );
   NAND2X1 i_21039 ( .Y (n_818),
	.B (n_796),
	.A (phi_6) );
   NAND2BX1 i_11 ( .Y (n_820),
	.B (ir[13]),
	.AN (ir[15]) );
   NOR2X1 i_1753 ( .Y (n_821),
	.B (n_820),
	.A (ir[14]) );
   NOR3X1 i_1750 ( .Y (n_823),
	.C (ir[14]),
	.B (ir[13]),
	.A (ir[15]) );
   NAND2X1 i_128 ( .Y (n_824),
	.B (n_4078),
	.A (ir[14]) );
   NAND2X1 i_3 ( .Y (n_828),
	.B (n_816),
	.A (n_793) );
   NAND2X1 i_21014 ( .Y (n_829),
	.B (n_783),
	.A (phi_3) );
   NAND3X1 i_174 ( .Y (n_830),
	.C (n_796),
	.B (n_794),
	.A (phi_6) );
   NAND2X1 i_153 ( .Y (n_831),
	.B (n_783),
	.A (phi_5) );
   NAND2X1 i_282 ( .Y (n_832),
	.B (n_4088),
	.A (ir[12]) );
   NOR2BX1 i_1702 ( .Y (n_835),
	.B (n_786),
	.AN (ir[12]) );
   AND2X1 i_77 ( .Y (n_836),
	.B (n_4087),
	.A (n_835) );
   NAND2X1 i_31 ( .Y (n_837),
	.B (ir[8]),
	.A (n_799) );
   NOR2BX1 i_172 ( .Y (n_838),
	.B (n_837),
	.AN (ir[11]) );
   AND2X1 i_207 ( .Y (n_839),
	.B (n_838),
	.A (n_835) );
   NAND2X1 i_26 ( .Y (n_840),
	.B (ir[11]),
	.A (ir[9]) );
   NOR2X1 i_33 ( .Y (n_841),
	.B (ir[8]),
	.A (ir[10]) );
   NAND2X1 i_171 ( .Y (n_842),
	.B (n_4085),
	.A (n_841) );
   NOR2X1 i_43 ( .Y (n_843),
	.B (n_4100),
	.A (ir[10]) );
   NOR2X1 i_50 ( .Y (n_844),
	.B (n_840),
	.A (n_788) );
   NOR4BX1 i_293 ( .Y (n_847),
	.D (n_4084),
	.C (n_844),
	.B (n_812),
	.AN (n_406) );
   NOR3X1 i_186 ( .Y (n_850),
	.C (n_818),
	.B (n_786),
	.A (ir[12]) );
   NAND2X1 i_188 ( .Y (n_851),
	.B (n_850),
	.A (n_794) );
   OAI21XL i_80 ( .Y (n_855),
	.B0 (n_813),
	.A1 (n_816),
	.A0 (ir[12]) );
   NOR2BX1 i_318 ( .Y (n_856),
	.B (update_stall),
	.AN (update_it) );
   NAND4X1 i_39 ( .Y (n_859),
	.D (n_4220),
	.C (n_856),
	.B (phi_6),
	.A (ir[7]) );
   NAND3X1 i_1937 ( .Y (n_863),
	.C (n_4078),
	.B (ir[12]),
	.A (ir[14]) );
   NAND2BX1 i_2207 ( .Y (n_864),
	.B (n_844),
	.AN (n_863) );
   NOR2BX1 i_187 ( .Y (n_865),
	.B (ir[6]),
	.AN (ir[7]) );
   NAND4BXL i_40 ( .Y (n_868),
	.D (n_865),
	.C (n_478),
	.B (ir[3]),
	.AN (n_864) );
   NOR2BX1 i_206 ( .Y (n_869),
	.B (n_868),
	.AN (ir[1]) );
   NOR2X1 i_1935 ( .Y (n_871),
	.B (ir[12]),
	.A (n_824) );
   NAND2X1 i_41 ( .Y (n_872),
	.B (n_791),
	.A (n_871) );
   NOR2X1 i_127 ( .Y (n_873),
	.B (n_864),
	.A (ir[0]) );
   NOR4X1 i_162 ( .Y (n_875),
	.D (ir[2]),
	.C (ir[1]),
	.B (n_864),
	.A (ir[0]) );
   NOR2BX1 i_205 ( .Y (n_876),
	.B (ir[5]),
	.AN (ir[4]) );
   NOR2BX1 i_333 ( .Y (n_877),
	.B (ir[3]),
	.AN (n_865) );
   AOI33X1 i_7 ( .Y (n_879),
	.B2 (n_791),
	.B1 (n_841),
	.B0 (n_871),
	.A2 (n_875),
	.A1 (n_877),
	.A0 (n_876) );
   NAND2X1 i_60 ( .Y (n_880),
	.B (n_879),
	.A (n_380) );
   AOI31X1 i_75 ( .Y (n_882),
	.B0 (n_880),
	.A2 (n_4082),
	.A1 (n_4092),
	.A0 (three_cycle) );
   AOI21X1 i_17 ( .Y (n_883),
	.B0 (n_704),
	.A1 (n_801),
	.A0 (n_871) );
   NOR2X1 i_160 ( .Y (n_884),
	.B (ir[9]),
	.A (ir[11]) );
   AOI32X1 i_8 ( .Y (n_886),
	.B1 (n_810),
	.B0 (n_841),
	.A2 (n_4087),
	.A1 (n_809),
	.A0 (n_884) );
   NOR2X1 i_47 ( .Y (n_889),
	.B (n_837),
	.A (ir[11]) );
   NAND2X1 i_2132 ( .Y (n_890),
	.B (n_871),
	.A (n_889) );
   NOR2X1 i_201 ( .Y (n_893),
	.B (n_806),
	.A (n_840) );
   NOR2X1 i_350 ( .Y (n_895),
	.B (skip_one),
	.A (two_cycle) );
   NAND2X1 i_21079 ( .Y (n_896),
	.B (n_895),
	.A (phi_6) );
   NOR2BX1 i_363 ( .Y (n_897),
	.B (ir[9]),
	.AN (gz) );
   AOI222X1 i_365 ( .Y (n_899),
	.C1 (n_4085),
	.C0 (nz),
	.B1 (n_884),
	.B0 (arnz),
	.A1 (n_897),
	.A0 (ir[11]) );
   NAND3BX1 i_357 ( .Y (n_902),
	.C (n_432),
	.B (n_431),
	.AN (n_812) );
   NAND3X1 i_376 ( .Y (n_905),
	.C (three_cycle),
	.B (n_794),
	.A (phi_6) );
   NOR2BX1 i_204 ( .Y (n_908),
	.B (ir[4]),
	.AN (ir[5]) );
   NOR2X1 i_46 ( .Y (n_910),
	.B (phi_1),
	.A (n_1105) );
   AOI22X1 i_1987 ( .Y (n_912),
	.B1 (n_4100),
	.B0 (n_4086),
	.A1 (n_871),
	.A0 (n_455) );
   NAND2BX1 i_36 ( .Y (n_913),
	.B (ir[11]),
	.AN (n_863) );
   AOI21X1 i_393 ( .Y (n_914),
	.B0 (n_823),
	.A1 (n_808),
	.A0 (ir[12]) );
   OAI21XL i_394 ( .Y (n_915),
	.B0 (n_914),
	.A1 (n_804),
	.A0 (n_4092) );
   AOI211X1 i_396 ( .Y (n_917),
	.C0 (n_483),
	.B0 (n_915),
	.A1 (n_836),
	.A0 (n_884) );
   NOR3X1 i_6 ( .Y (n_920),
	.C (n_820),
	.B (n_1105),
	.A (ir[14]) );
   NAND2X1 i_4 ( .Y (n_922),
	.B (n_4221),
	.A (n_794) );
   NOR2X1 i_192 ( .Y (n_923),
	.B (n_818),
	.A (n_922) );
   NAND2X1 i_51 ( .Y (n_924),
	.B (n_4076),
	.A (phi_6) );
   NAND2BX1 i_18 ( .Y (n_925),
	.B (n_382),
	.AN (n_467) );
   NAND2X1 i_1858 ( .Y (n_926),
	.B (n_810),
	.A (n_843) );
   NAND2X1 i_118 ( .Y (n_927),
	.B (n_886),
	.A (n_926) );
   AOI211X1 i_406 ( .Y (n_928),
	.C0 (ir[14]),
	.B0 (ir[15]),
	.A1 (ir[12]),
	.A0 (ir[13]) );
   NOR3X1 i_81 ( .Y (n_930),
	.C (n_925),
	.B (n_928),
	.A (n_927) );
   NAND2X1 i_61 ( .Y (n_931),
	.B (n_883),
	.A (n_890) );
   OAI21XL i_9 ( .Y (n_932),
	.B0 (n_4091),
	.A1 (n_913),
	.A0 (n_837) );
   AOI32X1 i_72 ( .Y (n_934),
	.B1 (n_812),
	.B0 (n_871),
	.A2 (n_869),
	.A1 (n_873),
	.A0 (ir[2]) );
   NOR2BX1 i_2194 ( .Y (n_935),
	.B (n_863),
	.AN (n_893) );
   AOI21X1 i_119 ( .Y (n_936),
	.B0 (n_935),
	.A1 (n_4087),
	.A0 (n_4086) );
   NAND2X1 i_19 ( .Y (n_937),
	.B (n_936),
	.A (n_934) );
   NOR4BX1 i_113 ( .Y (n_940),
	.D (n_931),
	.C (n_932),
	.B (n_937),
	.AN (n_930) );
   NOR3X1 i_49 ( .Y (n_941),
	.C (reset),
	.B (phi_1),
	.A (n_1105) );
   AOI22X1 i_82 ( .Y (n_943),
	.B1 (n_802),
	.B0 (ir[12]),
	.A1 (n_787),
	.A0 (n_793) );
   AOI221XL i_430 ( .Y (n_945),
	.C0 (n_584),
	.B1 (n_836),
	.B0 (ir[9]),
	.A1 (n_485),
	.A0 (n_835) );
   NOR2X1 i_114 ( .Y (n_948),
	.B (reset),
	.A (n_859) );
   NOR2BX1 i_435 ( .Y (n_949),
	.B (n_493),
	.AN (n_1105) );
   NOR2BX1 i_138 ( .Y (n_950),
	.B (n_932),
	.AN (n_382) );
   NAND2X1 i_184 ( .Y (n_951),
	.B (n_864),
	.A (n_950) );
   NOR3X1 i_2136 ( .Y (n_952),
	.C (n_790),
	.B (ir[12]),
	.A (n_824) );
   SDFFRHQX1 branch_stall_delay_reg ( .SI (BG_scan_in),
	.SE (scan_en),
	.RN (n_4221),
	.Q (branch_stall_delay),
	.D (n_3104),
	.CK (clk) );
   OAI21XL i_3342 ( .Y (n_3104),
	.B0 (n_3107),
	.A1 (n_1103),
	.A0 (n_2515) );
   NAND2X1 i_3344 ( .Y (n_3107),
	.B (branch_stall_delay),
	.A (n_2515) );
   NOR2X1 i_139 ( .Y (n_954),
	.B (n_952),
	.A (n_496) );
   SDFFRHQX1 branch_stall_reg ( .SI (branch_stall_delay),
	.SE (FE_OFN163_scan_enI),
	.RN (n_4221),
	.Q (branch_stall),
	.D (n_3110),
	.CK (clk) );
   OAI31X1 i_3349 ( .Y (n_3110),
	.B0 (n_3113),
	.A2 (n_4083),
	.A1 (n_407),
	.A0 (n_383) );
   NAND3X1 i_3352 ( .Y (n_3113),
	.C (n_1103),
	.B (branch_stall),
	.A (n_407) );
   NAND2BX1 i_442 ( .Y (n_955),
	.B (n_890),
	.AN (n_704) );
   SDFFRHQX1 update_stall_reg ( .SI (branch_stall),
	.SE (scan_en),
	.RN (n_4221),
	.Q (update_stall),
	.D (n_3116),
	.CK (clk) );
   MX2X1 i_3357 ( .Y (n_3116),
	.S0 (phi_1),
	.B (branch_stall),
	.A (update_stall) );
   SDFFRHQX1 three_cycle_reg ( .SI (update_stall),
	.SE (FE_OFN165_scan_enI),
	.RN (n_4221),
	.Q (three_cycle),
	.D (n_3122),
	.CK (clk) );
   MX2X1 i_3364 ( .Y (n_3122),
	.S0 (n_2765),
	.B (n_2768),
	.A (three_cycle) );
   SDFFRHQX1 two_cycle_reg ( .SI (three_cycle),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (two_cycle),
	.D (n_4093),
	.CK (clk) );
   AOI21X1 i_3371 ( .Y (n_3128),
	.B0 (n_3130),
	.A1 (two_cycle),
	.A0 (n_1833) );
   AOI31X1 i_3372 ( .Y (n_3130),
	.B0 (n_1833),
	.A2 (n_1111),
	.A1 (n_1062),
	.A0 (n_1114) );
   SDFFRHQX1 update_it_reg ( .SI (two_cycle),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (update_it),
	.D (n_3134),
	.CK (clk) );
   OAI21XL i_3378 ( .Y (n_3134),
	.B0 (n_3137),
	.A1 (n_3146),
	.A0 (n_1105) );
   NAND2X1 i_3380 ( .Y (n_3137),
	.B (update_it),
	.A (n_3146) );
   NAND2X1 i_48 ( .Y (n_959),
	.B (n_4076),
	.A (phi_3) );
   SDFFHQX1 acc_reg_0 ( .SI (update_it),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[0]),
	.D (n_3140),
	.CK (clk) );
   OAI2BB1X1 i_3385 ( .Y (n_3140),
	.B0 (n_3142),
	.A1N (acc[0]),
	.A0N (n_4094) );
   NAND2X1 i_3386 ( .Y (n_3142),
	.B (\nbus_440[0] ),
	.A (alu_result[0]) );
   NOR2X1 i_449 ( .Y (n_960),
	.B (n_4077),
	.A (n_959) );
   SEDFFX1 acc_reg_1 ( .SI (acc[0]),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[1]),
	.E (\nbus_440[0] ),
	.D (alu_result[1]),
	.CK (clk) );
   SEDFFX1 acc_reg_2 ( .SI (acc[1]),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[2]),
	.E (\nbus_440[0] ),
	.D (alu_result[2]),
	.CK (clk) );
   NOR2X1 i_135 ( .Y (n_962),
	.B (n_584),
	.A (n_952) );
   SEDFFX1 acc_reg_3 ( .SI (acc[2]),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[3]),
	.E (\nbus_440[0] ),
	.D (alu_result[3]),
	.CK (clk) );
   SEDFFX1 acc_reg_4 ( .SI (acc[3]),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[4]),
	.E (\nbus_440[0] ),
	.D (alu_result[4]),
	.CK (clk) );
   SEDFFX1 acc_reg_5 ( .SI (acc[4]),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[5]),
	.E (\nbus_440[0] ),
	.D (alu_result[5]),
	.CK (clk) );
   NAND2X1 i_140 ( .Y (n_965),
	.B (pc[14]),
	.A (pc[11]) );
   SEDFFX1 acc_reg_6 ( .SI (acc[5]),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[6]),
	.E (\nbus_440[0] ),
	.D (alu_result[6]),
	.CK (clk) );
   NAND2X1 i_1 ( .Y (n_966),
	.B (pc[1]),
	.A (pc[0]) );
   SEDFFX1 acc_reg_7 ( .SI (acc[6]),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[7]),
	.E (\nbus_440[0] ),
	.D (alu_result[7]),
	.CK (clk) );
   NAND3X1 i_58 ( .Y (n_967),
	.C (pc[2]),
	.B (pc[1]),
	.A (pc[0]) );
   SEDFFX1 acc_reg_8 ( .SI (acc[7]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[8]),
	.E (\nbus_440[0] ),
	.D (alu_result[8]),
	.CK (clk) );
   NAND2BX1 i_108 ( .Y (n_968),
	.B (pc[3]),
	.AN (n_967) );
   SEDFFX1 acc_reg_9 ( .SI (acc[8]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[9]),
	.E (\nbus_440[0] ),
	.D (alu_result[9]),
	.CK (clk) );
   NAND2BX1 i_361755 ( .Y (n_969),
	.B (pc[4]),
	.AN (n_968) );
   SEDFFX1 acc_reg_10 ( .SI (acc[9]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[10]),
	.E (\nbus_440[0] ),
	.D (alu_result[10]),
	.CK (clk) );
   NAND2BX1 i_56 ( .Y (n_970),
	.B (pc[5]),
	.AN (n_969) );
   SEDFFX1 acc_reg_11 ( .SI (acc[10]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[11]),
	.E (\nbus_440[0] ),
	.D (alu_result[11]),
	.CK (clk) );
   NAND2BX1 i_107 ( .Y (n_971),
	.B (pc[6]),
	.AN (n_970) );
   SEDFFX1 acc_reg_12 ( .SI (acc[11]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[12]),
	.E (\nbus_440[0] ),
	.D (alu_result[12]),
	.CK (clk) );
   NAND2BX1 i_30 ( .Y (n_972),
	.B (pc[7]),
	.AN (n_971) );
   SEDFFX1 acc_reg_13 ( .SI (acc[12]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[13]),
	.E (\nbus_440[0] ),
	.D (alu_result[13]),
	.CK (clk) );
   NAND2BX1 i_143 ( .Y (n_973),
	.B (pc[8]),
	.AN (n_972) );
   SEDFFX1 acc_reg_14 ( .SI (acc[13]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[14]),
	.E (\nbus_440[0] ),
	.D (alu_result[14]),
	.CK (clk) );
   NAND2BX1 i_57 ( .Y (n_974),
	.B (pc[9]),
	.AN (n_973) );
   SEDFFX1 acc_reg_15 ( .SI (acc[14]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[15]),
	.E (\nbus_440[0] ),
	.D (alu_result[15]),
	.CK (clk) );
   NAND2BX1 i_581765 ( .Y (n_975),
	.B (pc[10]),
	.AN (n_974) );
   SEDFFX1 acc_reg_16 ( .SI (acc[15]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[16]),
	.E (\nbus_440[0] ),
	.D (alu_result[16]),
	.CK (clk) );
   NAND2X1 i_68 ( .Y (n_976),
	.B (pc[12]),
	.A (pc[13]) );
   SEDFFX1 acc_reg_17 ( .SI (acc[16]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[17]),
	.E (\nbus_440[0] ),
	.D (alu_result[17]),
	.CK (clk) );
   SEDFFX1 acc_reg_18 ( .SI (acc[17]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[18]),
	.E (\nbus_440[0] ),
	.D (alu_result[18]),
	.CK (clk) );
   NOR3X1 i_159 ( .Y (n_978),
	.C (n_965),
	.B (n_976),
	.A (n_975) );
   SEDFFX1 acc_reg_19 ( .SI (acc[18]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[19]),
	.E (\nbus_440[0] ),
	.D (alu_result[19]),
	.CK (clk) );
   NAND2X1 i_42 ( .Y (n_979),
	.B (pc[11]),
	.A (pc[10]) );
   SEDFFX1 acc_reg_20 ( .SI (acc[19]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[20]),
	.E (\nbus_440[0] ),
	.D (alu_result[20]),
	.CK (clk) );
   SEDFFX1 acc_reg_21 ( .SI (acc[20]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[21]),
	.E (\nbus_440[0] ),
	.D (alu_result[21]),
	.CK (clk) );
   NOR3X1 i_156 ( .Y (n_981),
	.C (n_974),
	.B (n_976),
	.A (n_979) );
   SEDFFX1 acc_reg_22 ( .SI (acc[21]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[22]),
	.E (\nbus_440[0] ),
	.D (alu_result[22]),
	.CK (clk) );
   NAND3X1 i_69 ( .Y (n_982),
	.C (pc[9]),
	.B (pc[11]),
	.A (pc[10]) );
   SEDFFX1 acc_reg_23 ( .SI (acc[22]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[23]),
	.E (\nbus_440[0] ),
	.D (alu_result[23]),
	.CK (clk) );
   SEDFFX1 acc_reg_24 ( .SI (acc[23]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[24]),
	.E (\nbus_440[0] ),
	.D (alu_result[24]),
	.CK (clk) );
   NOR3X1 i_157 ( .Y (n_984),
	.C (n_4101),
	.B (n_982),
	.A (n_973) );
   SEDFFX1 acc_reg_25 ( .SI (acc[24]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[25]),
	.E (\nbus_440[0] ),
	.D (alu_result[25]),
	.CK (clk) );
   SEDFFX1 acc_reg_26 ( .SI (acc[25]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[26]),
	.E (\nbus_440[0] ),
	.D (alu_result[26]),
	.CK (clk) );
   SEDFFX1 acc_reg_27 ( .SI (acc[26]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[27]),
	.E (\nbus_440[0] ),
	.D (alu_result[27]),
	.CK (clk) );
   SEDFFX1 acc_reg_28 ( .SI (acc[27]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[28]),
	.E (\nbus_440[0] ),
	.D (alu_result[28]),
	.CK (clk) );
   SEDFFX1 acc_reg_29 ( .SI (acc[28]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[29]),
	.E (\nbus_440[0] ),
	.D (alu_result[29]),
	.CK (clk) );
   NAND3X1 i_155 ( .Y (n_989),
	.C (n_4080),
	.B (n_886),
	.A (n_926) );
   SEDFFX1 acc_reg_30 ( .SI (acc[29]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[30]),
	.E (\nbus_440[0] ),
	.D (alu_result[30]),
	.CK (clk) );
   SEDFFX1 acc_reg_31 ( .SI (acc[30]),
	.SE (FE_OFN14_scan_enI),
	.Q (acc[31]),
	.E (\nbus_440[0] ),
	.D (alu_result[31]),
	.CK (clk) );
   SEDFFX1 acc_reg_32 ( .SI (acc[31]),
	.SE (FE_OFN9_scan_enI),
	.Q (acc[32]),
	.E (\nbus_440[0] ),
	.D (alu_result[32]),
	.CK (clk) );
   NAND3BX1 i_13 ( .Y (n_992),
	.C (n_1105),
	.B (n_876),
	.AN (arp) );
   SDFFRHQX1 arp_reg ( .SI (acc[32]),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (FE_OFN131_arp),
	.D (n_3340),
	.CK (clk) );
   OAI2BB1X1 i_3621 ( .Y (n_3340),
	.B0 (n_3343),
	.A1N (n_1104),
	.A0N (ir[0]) );
   NAND2BX1 i_3623 ( .Y (n_3343),
	.B (arp),
	.AN (n_1104) );
   SDFFHQX1 null_op_reg0 ( .SI (arp),
	.SE (FE_OFN139_scan_enI),
	.Q (Q),
	.D (n_3349),
	.CK (clk) );
   AND2X1 i_3630 ( .Y (n_3349),
	.B (Q),
	.A (n_2909) );
   OR3XL i_65 ( .Y (n_994),
	.C (ar[2]),
	.B (ar[1]),
	.A (ar[0]) );
   SDFFRHQX1 ovm_reg ( .SI (Q),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (ovm),
	.D (n_3352),
	.CK (clk) );
   OAI21XL i_3635 ( .Y (n_3352),
	.B0 (n_3354),
	.A1 (n_4223),
	.A0 (n_1108) );
   NAND4BXL i_3636 ( .Y (n_3354),
	.D (n_869),
	.C (n_1108),
	.B (ir[0]),
	.AN (ir[2]) );
   NOR2X1 i_98 ( .Y (n_995),
	.B (ar[3]),
	.A (n_994) );
   SEDFFX1 sel_op_b_reg_0 ( .SI (ovm),
	.SE (FE_OFN9_scan_enI),
	.Q (sel_op_b[0]),
	.E (\nbus_434[0] ),
	.D (nbus_439[0]),
	.CK (clk) );
   NOR2X1 i_129 ( .Y (n_996),
	.B (ar[4]),
	.A (n_4074) );
   SEDFFX1 sel_op_b_reg_1 ( .SI (sel_op_b[0]),
	.SE (FE_OFN9_scan_enI),
	.Q (sel_op_b[1]),
	.E (\nbus_434[0] ),
	.D (nbus_439[1]),
	.CK (clk) );
   OR3XL i_130 ( .Y (n_997),
	.C (n_4074),
	.B (ar[5]),
	.A (ar[4]) );
   SEDFFX1 sel_op_b_reg_2 ( .SI (sel_op_b[1]),
	.SE (FE_OFN9_scan_enI),
	.Q (sel_op_b[2]),
	.E (\nbus_434[0] ),
	.D (nbus_439[2]),
	.CK (clk) );
   NOR2X1 i_131 ( .Y (n_998),
	.B (ar[6]),
	.A (n_997) );
   SDFFRHQX1 skip_one_reg ( .SI (sel_op_b[2]),
	.SE (scan_en),
	.RN (n_4221),
	.Q (skip_one),
	.D (n_3376),
	.CK (clk) );
   OAI21XL i_3664 ( .Y (n_3376),
	.B0 (n_3379),
	.A1 (n_1790),
	.A0 (n_1793) );
   NAND2X1 i_3666 ( .Y (n_3379),
	.B (skip_one),
	.A (n_1790) );
   NOR2X1 i_34 ( .Y (n_999),
	.B (ar[7]),
	.A (n_4073) );
   SDFFRHQX1 ov_flag_reg ( .SI (skip_one),
	.SE (FE_OFN163_scan_enI),
	.RN (n_4221),
	.Q (ov),
	.D (n_3382),
	.CK (clk) );
   OAI21XL i_3671 ( .Y (n_3382),
	.B0 (n_3385),
	.A1 (n_2384),
	.A0 (n_2387) );
   NAND2X1 i_3673 ( .Y (n_3385),
	.B (ov),
	.A (n_2384) );
   OR3XL i_163 ( .Y (n_1000),
	.C (n_4073),
	.B (ar[8]),
	.A (ar[7]) );
   SDFFSHQX1 pc_reg_0 ( .SN (n_4221),
	.SI (ov),
	.SE (FE_OFN163_scan_enI),
	.Q (pc[0]),
	.D (n_3388),
	.CK (clk) );
   MX2X1 i_3678 ( .Y (n_3388),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[0]),
	.A (pc[0]) );
   NOR2X1 i_164 ( .Y (n_1001),
	.B (ar[9]),
	.A (n_1000) );
   SDFFSHQX1 pc_reg_1 ( .SN (n_4221),
	.SI (pc[0]),
	.SE (scan_en),
	.Q (pc[1]),
	.D (n_3394),
	.CK (clk) );
   MX2X1 i_3685 ( .Y (n_3394),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[1]),
	.A (pc[1]) );
   NOR2X1 i_165 ( .Y (n_1002),
	.B (ar[10]),
	.A (n_4072) );
   SDFFSHQX1 pc_reg_2 ( .SN (n_4221),
	.SI (pc[1]),
	.SE (scan_en),
	.Q (pc[2]),
	.D (n_3400),
	.CK (clk) );
   MX2X1 i_3692 ( .Y (n_3400),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[2]),
	.A (pc[2]) );
   SDFFSHQX1 pc_reg_3 ( .SN (n_4221),
	.SI (pc[2]),
	.SE (scan_en),
	.Q (pc[3]),
	.D (n_3406),
	.CK (clk) );
   MX2X1 i_3699 ( .Y (n_3406),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[3]),
	.A (pc[3]) );
   SDFFSHQX1 pc_reg_4 ( .SN (n_4221),
	.SI (pc[3]),
	.SE (FE_OFN166_scan_enI),
	.Q (pc[4]),
	.D (n_3412),
	.CK (clk) );
   MX2X1 i_3706 ( .Y (n_3412),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[4]),
	.A (pc[4]) );
   NOR4X1 i_566 ( .Y (n_1005),
	.D (ar[14]),
	.C (ar[13]),
	.B (ar[12]),
	.A (ar[11]) );
   SDFFSHQX1 pc_reg_5 ( .SN (n_4221),
	.SI (pc[4]),
	.SE (FE_OFN166_scan_enI),
	.Q (pc[5]),
	.D (n_3418),
	.CK (clk) );
   MX2X1 i_3713 ( .Y (n_3418),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[5]),
	.A (pc[5]) );
   NAND2X1 i_169 ( .Y (n_1006),
	.B (n_1005),
	.A (n_1002) );
   SDFFSHQX1 pc_reg_6 ( .SN (n_4221),
	.SI (pc[5]),
	.SE (FE_OFN164_scan_enI),
	.Q (pc[6]),
	.D (n_3424),
	.CK (clk) );
   MX2X1 i_3720 ( .Y (n_3424),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[6]),
	.A (pc[6]) );
   SDFFSHQX1 pc_reg_7 ( .SN (n_4221),
	.SI (pc[6]),
	.SE (FE_OFN164_scan_enI),
	.Q (pc[7]),
	.D (n_3430),
	.CK (clk) );
   MX2X1 i_3727 ( .Y (n_3430),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[7]),
	.A (pc[7]) );
   NAND3BX1 i_12 ( .Y (n_1008),
	.C (n_1105),
	.B (n_908),
	.AN (arp) );
   SDFFSHQX1 pc_reg_8 ( .SN (n_4221),
	.SI (pc[7]),
	.SE (scan_en),
	.Q (pc[8]),
	.D (n_3436),
	.CK (clk) );
   MX2X1 i_3735 ( .Y (n_3436),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[8]),
	.A (pc[8]) );
   NAND2X1 i_12042 ( .Y (n_1009),
	.B (ar[1]),
	.A (ar[0]) );
   SDFFSHQX1 pc_reg_9 ( .SN (n_4221),
	.SI (pc[8]),
	.SE (scan_en),
	.Q (pc[9]),
	.D (n_3442),
	.CK (clk) );
   MX2X1 i_3743 ( .Y (n_3442),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[9]),
	.A (pc[9]) );
   NAND3X1 i_64 ( .Y (n_1010),
	.C (ar[2]),
	.B (ar[1]),
	.A (ar[0]) );
   SDFFSHQX1 pc_reg_10 ( .SN (n_4221),
	.SI (pc[9]),
	.SE (FE_OFN162_scan_enI),
	.Q (pc[10]),
	.D (n_3448),
	.CK (clk) );
   MX2X1 i_3751 ( .Y (n_3448),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[10]),
	.A (pc[10]) );
   NAND2BX1 i_192059 ( .Y (n_1011),
	.B (ar[3]),
	.AN (n_1010) );
   SDFFSHQX1 pc_reg_11 ( .SN (n_4221),
	.SI (pc[10]),
	.SE (FE_OFN162_scan_enI),
	.Q (pc[11]),
	.D (n_3454),
	.CK (clk) );
   MX2X1 i_3758 ( .Y (n_3454),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[11]),
	.A (pc[11]) );
   NAND2BX1 i_59 ( .Y (n_1012),
	.B (ar[4]),
	.AN (n_1011) );
   SDFFSHQX1 pc_reg_12 ( .SN (n_4221),
	.SI (pc[11]),
	.SE (scan_en),
	.Q (pc[12]),
	.D (n_3460),
	.CK (clk) );
   MXI2X1 i_3765 ( .Y (n_3460),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[12]),
	.A (n_4101) );
   NAND2BX1 i_372075 ( .Y (n_1013),
	.B (ar[5]),
	.AN (n_1012) );
   SDFFSHQX1 pc_reg_13 ( .SN (n_4221),
	.SI (pc[12]),
	.SE (FE_OFN162_scan_enI),
	.Q (pc[13]),
	.D (n_3466),
	.CK (clk) );
   MX2X1 i_3772 ( .Y (n_3466),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[13]),
	.A (pc[13]) );
   NAND2BX1 i_382076 ( .Y (n_1014),
	.B (ar[6]),
	.AN (n_1013) );
   SDFFSHQX1 pc_reg_14 ( .SN (n_4221),
	.SI (pc[13]),
	.SE (scan_en),
	.Q (pc[14]),
	.D (n_3472),
	.CK (clk) );
   MX2X1 i_3779 ( .Y (n_3472),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[14]),
	.A (pc[14]) );
   NAND2BX1 i_53 ( .Y (n_1015),
	.B (ar[7]),
	.AN (n_1014) );
   SDFFSHQX1 pc_reg_15 ( .SN (n_4221),
	.SI (pc[14]),
	.SE (scan_en),
	.Q (pc[15]),
	.D (n_3478),
	.CK (clk) );
   MX2X1 i_3786 ( .Y (n_3478),
	.S0 (\nbus_436[0] ),
	.B (nbus_437[15]),
	.A (pc[15]) );
   SDFFRHQX1 read_prog_reg ( .SI (pc[15]),
	.SE (scan_en),
	.RN (n_4221),
	.Q (read_prog),
	.D (n_3484),
	.CK (clk) );
   OAI21XL i_3793 ( .Y (n_3484),
	.B0 (n_3487),
	.A1 (n_1940),
	.A0 (n_2610) );
   NAND2X1 i_3795 ( .Y (n_3487),
	.B (read_prog),
	.A (n_1940) );
   NAND3BX1 i_191 ( .Y (n_1017),
	.C (ar[8]),
	.B (ar[9]),
	.AN (n_1015) );
   SDFFRHQX1 dp_reg ( .SI (read_prog),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (dp),
	.D (n_3490),
	.CK (clk) );
   OAI21XL i_3800 ( .Y (n_3490),
	.B0 (n_3493),
	.A1 (n_1107),
	.A0 (n_2534) );
   NAND2X1 i_3802 ( .Y (n_3493),
	.B (dp),
	.A (n_1107) );
   NAND2BX1 i_582093 ( .Y (n_1018),
	.B (ar[10]),
	.AN (n_1017) );
   SEDFFX1 sel_op_a_reg_0 ( .SI (dp),
	.SE (FE_OFN9_scan_enI),
	.Q (sel_op_a[0]),
	.E (\nbus_434[0] ),
	.D (nbus_435[0]),
	.CK (clk) );
   SEDFFX1 sel_op_a_reg_1 ( .SI (sel_op_a[0]),
	.SE (FE_OFN9_scan_enI),
	.Q (sel_op_a[1]),
	.E (\nbus_434[0] ),
	.D (nbus_435[1]),
	.CK (clk) );
   SEDFFX1 sel_op_a_reg_2 ( .SI (sel_op_a[1]),
	.SE (FE_OFN9_scan_enI),
	.Q (sel_op_a[2]),
	.E (\nbus_434[0] ),
	.D (nbus_435[2]),
	.CK (clk) );
   NAND4X1 i_561 ( .Y (n_1021),
	.D (ar[13]),
	.C (ar[14]),
	.B (ar[12]),
	.A (ar[11]) );
   SDFFRHQX1 go_port_reg ( .SI (sel_op_a[2]),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (go_port),
	.D (n_3514),
	.CK (clk) );
   OAI31X1 i_3828 ( .Y (n_3514),
	.B0 (n_3517),
	.A2 (n_832),
	.A1 (n_2115),
	.A0 (n_830) );
   NAND2X1 i_3830 ( .Y (n_3517),
	.B (go_port),
	.A (n_2115) );
   NOR2X1 i_622097 ( .Y (n_1022),
	.B (n_1021),
	.A (n_1018) );
   SEDFFX1 top_reg_0 ( .SI (go_port),
	.SE (scan_en),
	.Q (top[0]),
	.E (\nbus_432[0] ),
	.D (mdr[0]),
	.CK (clk) );
   SEDFFX1 top_reg_1 ( .SI (top[0]),
	.SE (scan_en),
	.Q (top[1]),
	.E (\nbus_432[0] ),
	.D (mdr[1]),
	.CK (clk) );
   SEDFFX1 top_reg_2 ( .SI (top[1]),
	.SE (scan_en),
	.Q (top[2]),
	.E (\nbus_432[0] ),
	.D (mdr[2]),
	.CK (clk) );
   OR3XL i_166 ( .Y (n_1025),
	.C (n_4072),
	.B (ar[11]),
	.A (ar[10]) );
   SEDFFX1 top_reg_3 ( .SI (top[2]),
	.SE (scan_en),
	.Q (top[3]),
	.E (\nbus_432[0] ),
	.D (mdr[3]),
	.CK (clk) );
   NOR2X1 i_167 ( .Y (n_1026),
	.B (n_1025),
	.A (ar[12]) );
   SEDFFX1 top_reg_4 ( .SI (top[3]),
	.SE (scan_en),
	.Q (top[4]),
	.E (\nbus_432[0] ),
	.D (mdr[4]),
	.CK (clk) );
   NOR2X1 i_168 ( .Y (n_1027),
	.B (ar[13]),
	.A (n_4075) );
   SEDFFX1 top_reg_5 ( .SI (top[4]),
	.SE (scan_en),
	.Q (top[5]),
	.E (\nbus_432[0] ),
	.D (mdr[5]),
	.CK (clk) );
   NAND2X1 i_197 ( .Y (n_1028),
	.B (ar[10]),
	.A (ar[11]) );
   SEDFFX1 top_reg_6 ( .SI (top[5]),
	.SE (scan_en),
	.Q (top[6]),
	.E (\nbus_432[0] ),
	.D (mdr[6]),
	.CK (clk) );
   NOR2X1 i_592094 ( .Y (n_1029),
	.B (n_1028),
	.A (n_1017) );
   SEDFFX1 top_reg_7 ( .SI (top[6]),
	.SE (scan_en),
	.Q (top[7]),
	.E (\nbus_432[0] ),
	.D (mdr[7]),
	.CK (clk) );
   SEDFFX1 top_reg_8 ( .SI (top[7]),
	.SE (scan_en),
	.Q (top[8]),
	.E (\nbus_432[0] ),
	.D (mdr[8]),
	.CK (clk) );
   NAND3X1 i_612096 ( .Y (n_1031),
	.C (n_1029),
	.B (ar[12]),
	.A (ar[13]) );
   SEDFFX1 top_reg_9 ( .SI (top[8]),
	.SE (scan_en),
	.Q (top[9]),
	.E (\nbus_432[0] ),
	.D (mdr[9]),
	.CK (clk) );
   SEDFFX1 top_reg_10 ( .SI (top[9]),
	.SE (scan_en),
	.Q (top[10]),
	.E (\nbus_432[0] ),
	.D (mdr[10]),
	.CK (clk) );
   NAND2BX1 i_562091 ( .Y (n_1033),
	.B (ar[8]),
	.AN (n_1015) );
   SEDFFX1 top_reg_11 ( .SI (top[10]),
	.SE (scan_en),
	.Q (top[11]),
	.E (\nbus_432[0] ),
	.D (mdr[11]),
	.CK (clk) );
   SEDFFX1 top_reg_12 ( .SI (top[11]),
	.SE (FE_OFN142_scan_enI),
	.Q (top[12]),
	.E (\nbus_432[0] ),
	.D (mdr[12]),
	.CK (clk) );
   NAND4X1 i_585 ( .Y (n_1035),
	.D (ar[9]),
	.C (ar[12]),
	.B (ar[10]),
	.A (ar[11]) );
   SEDFFX1 top_reg_13 ( .SI (top[12]),
	.SE (FE_OFN142_scan_enI),
	.Q (top[13]),
	.E (\nbus_432[0] ),
	.D (mdr[13]),
	.CK (clk) );
   OR2X1 i_602095 ( .Y (n_1036),
	.B (n_1035),
	.A (n_1033) );
   SEDFFX1 top_reg_14 ( .SI (top[13]),
	.SE (scan_en),
	.Q (top[14]),
	.E (\nbus_432[0] ),
	.D (mdr[14]),
	.CK (clk) );
   SEDFFX1 top_reg_15 ( .SI (top[14]),
	.SE (scan_en),
	.Q (top[15]),
	.E (\nbus_432[0] ),
	.D (mdr[15]),
	.CK (clk) );
   SDFFRHQX1 dmov_inc_reg ( .SI (top[15]),
	.SE (scan_en),
	.RN (n_4221),
	.Q (FE_OFN129_dmov_inc),
	.D (n_3616),
	.CK (clk) );
   MX2X1 i_3949 ( .Y (n_3616),
	.S0 (n_2235),
	.B (n_4081),
	.A (dmov_inc) );
   SDFFRHQX1 read_data_reg ( .SI (dmov_inc),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (read_data),
	.D (n_3625),
	.CK (clk) );
   AND2X1 i_3958 ( .Y (n_3625),
	.B (read_data),
	.A (n_2079) );
   SDFFRHQX1 read_port_reg ( .SI (read_data),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (read_port),
	.D (n_3631),
	.CK (clk) );
   AND2X1 i_3966 ( .Y (n_3631),
	.B (read_port),
	.A (n_2115) );
   SDFFRHQX1 go_data_reg ( .SI (read_port),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (go_data),
	.D (n_3634),
	.CK (clk) );
   OAI21XL i_3971 ( .Y (n_3634),
	.B0 (n_3637),
	.A1 (n_2082),
	.A0 (n_2079) );
   NAND2X1 i_3973 ( .Y (n_3637),
	.B (go_data),
	.A (n_2079) );
   SEDFFX1 ar0_reg_0 ( .SI (go_data),
	.SE (FE_OFN139_scan_enI),
	.Q (ar0[0]),
	.E (\nbus_430[0] ),
	.D (nbus_431[0]),
	.CK (clk) );
   NOR2X1 i_16 ( .Y (n_1043),
	.B (n_824),
	.A (n_1105) );
   SEDFFX1 ar0_reg_1 ( .SI (ar0[0]),
	.SE (scan_en),
	.Q (ar0[1]),
	.E (\nbus_430[0] ),
	.D (nbus_431[1]),
	.CK (clk) );
   AOI22X1 i_144 ( .Y (n_1044),
	.B1 (n_920),
	.B0 (mdr[7]),
	.A1 (n_1043),
	.A0 (ir[7]) );
   SEDFFX1 ar0_reg_2 ( .SI (ar0[1]),
	.SE (FE_OFN139_scan_enI),
	.Q (ar0[2]),
	.E (\nbus_430[0] ),
	.D (nbus_431[2]),
	.CK (clk) );
   AOI2BB1X1 i_642 ( .Y (n_1045),
	.B0 (n_644),
	.A1N (n_992),
	.A0N (n_751) );
   SEDFFX1 ar0_reg_3 ( .SI (ar0[2]),
	.SE (scan_en),
	.Q (ar0[3]),
	.E (\nbus_430[0] ),
	.D (nbus_431[3]),
	.CK (clk) );
   AOI22X1 i_145 ( .Y (n_1046),
	.B1 (n_920),
	.B0 (mdr[6]),
	.A1 (n_1043),
	.A0 (ir[6]) );
   SEDFFX1 ar0_reg_4 ( .SI (ar0[3]),
	.SE (scan_en),
	.Q (ar0[4]),
	.E (\nbus_430[0] ),
	.D (nbus_431[4]),
	.CK (clk) );
   AOI2BB1X1 i_651 ( .Y (n_1047),
	.B0 (n_651),
	.A1N (n_992),
	.A0N (n_755) );
   SEDFFX1 ar0_reg_5 ( .SI (ar0[4]),
	.SE (scan_en),
	.Q (ar0[5]),
	.E (\nbus_430[0] ),
	.D (nbus_431[5]),
	.CK (clk) );
   AOI22X1 i_146 ( .Y (n_1048),
	.B1 (n_920),
	.B0 (mdr[5]),
	.A1 (n_1043),
	.A0 (ir[5]) );
   SEDFFX1 ar0_reg_6 ( .SI (ar0[5]),
	.SE (scan_en),
	.Q (ar0[6]),
	.E (\nbus_430[0] ),
	.D (nbus_431[6]),
	.CK (clk) );
   AOI2BB1X1 i_660 ( .Y (n_1049),
	.B0 (n_658),
	.A1N (n_1008),
	.A0N (n_759) );
   SEDFFX1 ar0_reg_7 ( .SI (ar0[6]),
	.SE (FE_OFN13_scan_enI),
	.Q (ar0[7]),
	.E (\nbus_430[0] ),
	.D (nbus_431[7]),
	.CK (clk) );
   AOI22X1 i_147 ( .Y (n_1050),
	.B1 (n_920),
	.B0 (mdr[4]),
	.A1 (n_1043),
	.A0 (ir[4]) );
   SEDFFX1 ar0_reg_8 ( .SI (ar0[7]),
	.SE (scan_en),
	.Q (ar0[8]),
	.E (\nbus_430[0] ),
	.D (nbus_431[8]),
	.CK (clk) );
   AOI2BB1X1 i_669 ( .Y (n_1051),
	.B0 (n_665),
	.A1N (n_992),
	.A0N (n_763) );
   SEDFFX1 ar0_reg_9 ( .SI (ar0[8]),
	.SE (FE_OFN14_scan_enI),
	.Q (ar0[9]),
	.E (\nbus_430[0] ),
	.D (nbus_431[9]),
	.CK (clk) );
   AOI22X1 i_148 ( .Y (n_1052),
	.B1 (n_920),
	.B0 (mdr[3]),
	.A1 (n_1043),
	.A0 (ir[3]) );
   SEDFFX1 ar0_reg_10 ( .SI (ar0[9]),
	.SE (scan_en),
	.Q (ar0[10]),
	.E (\nbus_430[0] ),
	.D (nbus_431[10]),
	.CK (clk) );
   AOI2BB1X1 i_678 ( .Y (n_1053),
	.B0 (n_672),
	.A1N (n_992),
	.A0N (n_767) );
   SEDFFX1 ar0_reg_11 ( .SI (ar0[10]),
	.SE (scan_en),
	.Q (ar0[11]),
	.E (\nbus_430[0] ),
	.D (nbus_431[11]),
	.CK (clk) );
   AOI22X1 i_149 ( .Y (n_1054),
	.B1 (n_920),
	.B0 (mdr[2]),
	.A1 (n_1043),
	.A0 (ir[2]) );
   SEDFFX1 ar0_reg_12 ( .SI (ar0[11]),
	.SE (FE_OFN143_scan_enI),
	.Q (ar0[12]),
	.E (\nbus_430[0] ),
	.D (nbus_431[12]),
	.CK (clk) );
   AOI2BB1X1 i_687 ( .Y (n_1055),
	.B0 (n_679),
	.A1N (n_992),
	.A0N (n_771) );
   SEDFFX1 ar0_reg_13 ( .SI (ar0[12]),
	.SE (scan_en),
	.Q (ar0[13]),
	.E (\nbus_430[0] ),
	.D (nbus_431[13]),
	.CK (clk) );
   AOI22X1 i_150 ( .Y (n_1056),
	.B1 (n_920),
	.B0 (mdr[1]),
	.A1 (n_1043),
	.A0 (ir[1]) );
   SEDFFX1 ar0_reg_14 ( .SI (ar0[13]),
	.SE (scan_en),
	.Q (ar0[14]),
	.E (\nbus_430[0] ),
	.D (nbus_431[14]),
	.CK (clk) );
   OAI21XL i_105 ( .Y (n_1057),
	.B0 (n_1009),
	.A1 (ar[1]),
	.A0 (ar[0]) );
   SEDFFX1 ar0_reg_15 ( .SI (ar0[14]),
	.SE (scan_en),
	.Q (ar0[15]),
	.E (\nbus_430[0] ),
	.D (nbus_431[15]),
	.CK (clk) );
   MX2X1 i_693 ( .Y (n_1058),
	.S0 (n_1057),
	.B (n_992),
	.A (n_1008) );
   SDFFRHQX1 go_prog_reg ( .SI (ar0[15]),
	.SE (FE_OFN165_scan_enI),
	.RN (n_4221),
	.Q (go_prog),
	.D (n_3736),
	.CK (clk) );
   OAI21XL i_4092 ( .Y (n_3736),
	.B0 (n_3739),
	.A1 (n_1943),
	.A0 (n_1940) );
   NAND2X1 i_4094 ( .Y (n_3739),
	.B (go_prog),
	.A (n_1940) );
   SDFFRHQX1 fetch_branch_reg ( .SI (go_prog),
	.SE (scan_en),
	.RN (n_4221),
	.Q (fetch_branch),
	.D (n_4095),
	.CK (clk) );
   AOI31X1 i_4099 ( .Y (n_3742),
	.B0 (n_3744),
	.A2 (fetch_branch),
	.A1 (n_407),
	.A0 (n_1103) );
   AOI211X1 i_4100 ( .Y (n_3744),
	.C0 (n_407),
	.B0 (n_444),
	.A1 (branch_stall),
	.A0 (phi_1) );
   SDFFHQX1 alu_cmd_reg_0 ( .SI (fetch_branch),
	.SE (FE_OFN9_scan_enI),
	.Q (alu_cmd[0]),
	.D (n_4096),
	.CK (clk) );
   AOI21X1 i_4106 ( .Y (n_3748),
	.B0 (n_3750),
	.A1 (alu_cmd[0]),
	.A0 (\nbus_428[0] ) );
   AOI31X1 i_4107 ( .Y (n_3750),
	.B0 (\nbus_428[0] ),
	.A2 (n_1071),
	.A1 (n_879),
	.A0 (n_934) );
   AOI22X1 i_151 ( .Y (n_1061),
	.B1 (n_920),
	.B0 (mdr[0]),
	.A1 (n_1043),
	.A0 (ir[0]) );
   SDFFHQX1 alu_cmd_reg_1 ( .SI (alu_cmd[0]),
	.SE (FE_OFN14_scan_enI),
	.Q (alu_cmd[1]),
	.D (n_3754),
	.CK (clk) );
   OAI21XL i_4113 ( .Y (n_3754),
	.B0 (n_3757),
	.A1 (\nbus_429[1] ),
	.A0 (\nbus_428[0] ) );
   NAND2X1 i_4115 ( .Y (n_3757),
	.B (alu_cmd[1]),
	.A (\nbus_428[0] ) );
   AOI22X1 i_710 ( .Y (n_1062),
	.B1 (n_802),
	.B0 (n_829),
	.A1 (n_4088),
	.A0 (n_784) );
   SEDFFX1 alu_cmd_reg_2 ( .SI (alu_cmd[1]),
	.SE (FE_OFN14_scan_enI),
	.Q (alu_cmd[2]),
	.E (n_4097),
	.D (\nbus_429[2] ),
	.CK (clk) );
   SDFFHQX1 alu_cmd_reg_3 ( .SI (alu_cmd[2]),
	.SE (FE_OFN14_scan_enI),
	.Q (alu_cmd[3]),
	.D (n_3769),
	.CK (clk) );
   AND2X1 i_4129 ( .Y (n_3769),
	.B (\nbus_428[0] ),
	.A (alu_cmd[3]) );
   NAND2X1 i_714 ( .Y (n_1064),
	.B (n_817),
	.A (n_794) );
   SEDFFX1 p_reg_0 ( .SI (alu_cmd[3]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[0]),
	.E (\nbus_426[0] ),
	.D (mpy_result[0]),
	.CK (clk) );
   OAI21XL i_123 ( .Y (n_1065),
	.B0 (n_926),
	.A1 (n_820),
	.A0 (ir[14]) );
   SEDFFX1 p_reg_1 ( .SI (p[0]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[1]),
	.E (\nbus_426[0] ),
	.D (mpy_result[1]),
	.CK (clk) );
   SEDFFX1 p_reg_2 ( .SI (p[1]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[2]),
	.E (\nbus_426[0] ),
	.D (mpy_result[2]),
	.CK (clk) );
   SEDFFX1 p_reg_3 ( .SI (p[2]),
	.SE (scan_en),
	.Q (p[3]),
	.E (\nbus_426[0] ),
	.D (mpy_result[3]),
	.CK (clk) );
   AOI211X1 i_730 ( .Y (n_1068),
	.C0 (n_1065),
	.B0 (n_470),
	.A1 (n_823),
	.A0 (ir[12]) );
   SEDFFX1 p_reg_4 ( .SI (p[3]),
	.SE (scan_en),
	.Q (p[4]),
	.E (\nbus_426[0] ),
	.D (mpy_result[4]),
	.CK (clk) );
   SEDFFX1 p_reg_5 ( .SI (p[4]),
	.SE (scan_en),
	.Q (p[5]),
	.E (\nbus_426[0] ),
	.D (mpy_result[5]),
	.CK (clk) );
   SEDFFX1 p_reg_6 ( .SI (p[5]),
	.SE (scan_en),
	.Q (p[6]),
	.E (\nbus_426[0] ),
	.D (mpy_result[6]),
	.CK (clk) );
   NOR4BX1 i_733 ( .Y (n_1071),
	.D (n_705),
	.C (n_467),
	.B (n_704),
	.AN (n_1068) );
   SEDFFX1 p_reg_7 ( .SI (p[6]),
	.SE (scan_en),
	.Q (p[7]),
	.E (\nbus_426[0] ),
	.D (mpy_result[7]),
	.CK (clk) );
   SEDFFX1 p_reg_8 ( .SI (p[7]),
	.SE (scan_en),
	.Q (p[8]),
	.E (\nbus_426[0] ),
	.D (mpy_result[8]),
	.CK (clk) );
   SEDFFX1 p_reg_9 ( .SI (p[8]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[9]),
	.E (\nbus_426[0] ),
	.D (mpy_result[9]),
	.CK (clk) );
   SEDFFX1 p_reg_10 ( .SI (p[9]),
	.SE (FE_OFN146_scan_enI),
	.Q (p[10]),
	.E (\nbus_426[0] ),
	.D (mpy_result[10]),
	.CK (clk) );
   SEDFFX1 p_reg_11 ( .SI (p[10]),
	.SE (FE_OFN146_scan_enI),
	.Q (p[11]),
	.E (\nbus_426[0] ),
	.D (mpy_result[11]),
	.CK (clk) );
   NAND4BXL i_753 ( .Y (n_1076),
	.D (n_713),
	.C (n_790),
	.B (n_871),
	.AN (n_812) );
   SEDFFX1 p_reg_12 ( .SI (p[11]),
	.SE (FE_OFN146_scan_enI),
	.Q (p[12]),
	.E (\nbus_426[0] ),
	.D (mpy_result[12]),
	.CK (clk) );
   SEDFFX1 p_reg_13 ( .SI (p[12]),
	.SE (FE_OFN146_scan_enI),
	.Q (p[13]),
	.E (\nbus_426[0] ),
	.D (mpy_result[13]),
	.CK (clk) );
   SEDFFX1 p_reg_14 ( .SI (p[13]),
	.SE (scan_en),
	.Q (p[14]),
	.E (\nbus_426[0] ),
	.D (mpy_result[14]),
	.CK (clk) );
   SEDFFX1 p_reg_15 ( .SI (p[14]),
	.SE (FE_OFN145_scan_enI),
	.Q (p[15]),
	.E (\nbus_426[0] ),
	.D (mpy_result[15]),
	.CK (clk) );
   SEDFFX1 p_reg_16 ( .SI (p[15]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[16]),
	.E (\nbus_426[0] ),
	.D (mpy_result[16]),
	.CK (clk) );
   NAND4X1 i_756 ( .Y (n_1081),
	.D (n_716),
	.C (n_943),
	.B (n_714),
	.A (n_715) );
   SEDFFX1 p_reg_17 ( .SI (p[16]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[17]),
	.E (\nbus_426[0] ),
	.D (mpy_result[17]),
	.CK (clk) );
   SEDFFX1 p_reg_18 ( .SI (p[17]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[18]),
	.E (\nbus_426[0] ),
	.D (mpy_result[18]),
	.CK (clk) );
   SEDFFX1 p_reg_19 ( .SI (p[18]),
	.SE (FE_OFN145_scan_enI),
	.Q (p[19]),
	.E (\nbus_426[0] ),
	.D (mpy_result[19]),
	.CK (clk) );
   NAND3X1 i_159005 ( .Y (n_1084),
	.C (n_1105),
	.B (n_876),
	.A (arp) );
   SEDFFX1 p_reg_20 ( .SI (p[19]),
	.SE (scan_en),
	.Q (p[20]),
	.E (\nbus_426[0] ),
	.D (mpy_result[20]),
	.CK (clk) );
   SEDFFX1 p_reg_21 ( .SI (p[20]),
	.SE (FE_OFN171_scan_enI),
	.Q (p[21]),
	.E (\nbus_426[0] ),
	.D (mpy_result[21]),
	.CK (clk) );
   NAND3X1 i_14 ( .Y (n_1086),
	.C (n_908),
	.B (n_1105),
	.A (arp) );
   SEDFFX1 p_reg_22 ( .SI (p[21]),
	.SE (FE_OFN171_scan_enI),
	.Q (p[22]),
	.E (\nbus_426[0] ),
	.D (mpy_result[22]),
	.CK (clk) );
   SEDFFX1 p_reg_23 ( .SI (p[22]),
	.SE (scan_en),
	.Q (p[23]),
	.E (\nbus_426[0] ),
	.D (mpy_result[23]),
	.CK (clk) );
   SEDFFX1 p_reg_24 ( .SI (p[23]),
	.SE (scan_en),
	.Q (p[24]),
	.E (\nbus_426[0] ),
	.D (mpy_result[24]),
	.CK (clk) );
   SEDFFX1 p_reg_25 ( .SI (p[24]),
	.SE (scan_en),
	.Q (p[25]),
	.E (\nbus_426[0] ),
	.D (mpy_result[25]),
	.CK (clk) );
   SEDFFX1 p_reg_26 ( .SI (p[25]),
	.SE (scan_en),
	.Q (p[26]),
	.E (\nbus_426[0] ),
	.D (mpy_result[26]),
	.CK (clk) );
   SEDFFX1 p_reg_27 ( .SI (p[26]),
	.SE (scan_en),
	.Q (p[27]),
	.E (\nbus_426[0] ),
	.D (mpy_result[27]),
	.CK (clk) );
   SEDFFX1 p_reg_28 ( .SI (p[27]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[28]),
	.E (\nbus_426[0] ),
	.D (mpy_result[28]),
	.CK (clk) );
   SEDFFX1 p_reg_29 ( .SI (p[28]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[29]),
	.E (\nbus_426[0] ),
	.D (mpy_result[29]),
	.CK (clk) );
   SEDFFX1 p_reg_30 ( .SI (p[29]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[30]),
	.E (\nbus_426[0] ),
	.D (mpy_result[30]),
	.CK (clk) );
   SEDFFX1 p_reg_31 ( .SI (p[30]),
	.SE (FE_OFN17_scan_enI),
	.Q (p[31]),
	.E (\nbus_426[0] ),
	.D (mpy_result[31]),
	.CK (clk) );
   SDFFRHQX1 pc_acc_reg ( .SI (p[31]),
	.SE (FE_OFN9_scan_enI),
	.RN (n_4221),
	.Q (pc_acc),
	.D (n_3964),
	.CK (clk) );
   MXI2X1 i_4360 ( .Y (n_3964),
	.S0 (n_1439),
	.B (n_1114),
	.A (n_4222) );
   SDFFHQX1 null_op_reg ( .SI (pc_acc),
	.SE (FE_OFN9_scan_enI),
	.Q (Q175),
	.D (n_3973),
	.CK (clk) );
   AND2X1 i_4369 ( .Y (n_3973),
	.B (Q175),
	.A (n_1109) );
   SDFFHQX1 ar1_reg_0 ( .SI (Q175),
	.SE (FE_OFN9_scan_enI),
	.Q (ar1[0]),
	.D (n_4098),
	.CK (clk) );
   AOI21X1 i_4374 ( .Y (n_3976),
	.B0 (n_3978),
	.A1 (ar1[0]),
	.A0 (\nbus_424[0] ) );
   AOI21X1 i_4375 ( .Y (n_3978),
	.B0 (\nbus_424[0] ),
	.A1 (n_781),
	.A0 (n_1061) );
   SEDFFX1 ar1_reg_1 ( .SI (ar1[0]),
	.SE (scan_en),
	.Q (ar1[1]),
	.E (n_4099),
	.D (\nbus_425[1] ),
	.CK (clk) );
   SEDFFX1 ar1_reg_2 ( .SI (ar1[1]),
	.SE (scan_en),
	.Q (ar1[2]),
	.E (n_4099),
	.D (\nbus_425[2] ),
	.CK (clk) );
   SEDFFX1 ar1_reg_3 ( .SI (ar1[2]),
	.SE (scan_en),
	.Q (ar1[3]),
	.E (n_4099),
	.D (\nbus_425[3] ),
	.CK (clk) );
   SEDFFX1 ar1_reg_4 ( .SI (ar1[3]),
	.SE (scan_en),
	.Q (ar1[4]),
	.E (n_4099),
	.D (\nbus_425[4] ),
	.CK (clk) );
   NAND2X1 i_2 ( .Y (n_1103),
	.B (phi_1),
	.A (branch_stall) );
   SEDFFX1 ar1_reg_5 ( .SI (ar1[4]),
	.SE (FE_OFN13_scan_enI),
	.Q (ar1[5]),
	.E (n_4099),
	.D (\nbus_425[5] ),
	.CK (clk) );
   NOR3BX1 i_3521 ( .Y (n_1104),
	.C (ir[3]),
	.B (n_859),
	.AN (n_1105) );
   SEDFFX1 ar1_reg_6 ( .SI (ar1[5]),
	.SE (scan_en),
	.Q (ar1[6]),
	.E (n_4099),
	.D (\nbus_425[6] ),
	.CK (clk) );
   NAND2BX1 i_2925 ( .Y (n_1105),
	.B (phi_5),
	.AN (update_stall) );
   SEDFFX1 ar1_reg_7 ( .SI (ar1[6]),
	.SE (scan_en),
	.Q (ar1[7]),
	.E (n_4099),
	.D (\nbus_425[7] ),
	.CK (clk) );
   NOR2X1 i_2471 ( .Y (n_1106),
	.B (n_830),
	.A (n_832) );
   SEDFFX1 ar1_reg_8 ( .SI (ar1[7]),
	.SE (scan_en),
	.Q (ar1[8]),
	.E (n_4099),
	.D (\nbus_425[8] ),
	.CK (clk) );
   NAND4X1 i_3748 ( .Y (n_1107),
	.D (n_871),
	.C (n_429),
	.B (n_794),
	.A (phi_6) );
   SEDFFX1 ar1_reg_9 ( .SI (ar1[8]),
	.SE (scan_en),
	.Q (ar1[9]),
	.E (n_4099),
	.D (\nbus_425[9] ),
	.CK (clk) );
   AOI211X1 i_4043 ( .Y (n_1108),
	.C0 (branch_stall),
	.B0 (branch_stall_delay),
	.A1 (n_450),
	.A0 (n_1112) );
   SEDFFX1 ar1_reg_10 ( .SI (ar1[9]),
	.SE (scan_en),
	.Q (ar1[10]),
	.E (n_4099),
	.D (\nbus_425[10] ),
	.CK (clk) );
   OAI31X1 i_2860 ( .Y (n_1109),
	.B0 (n_4076),
	.A2 (n_712),
	.A1 (n_1081),
	.A0 (n_717) );
   SEDFFX1 ar1_reg_11 ( .SI (ar1[10]),
	.SE (scan_en),
	.Q (ar1[11]),
	.E (n_4099),
	.D (\nbus_425[11] ),
	.CK (clk) );
   SEDFFX1 ar1_reg_12 ( .SI (ar1[11]),
	.SE (FE_OFN143_scan_enI),
	.Q (ar1[12]),
	.E (n_4099),
	.D (\nbus_425[12] ),
	.CK (clk) );
   NAND2BX1 i_2475 ( .Y (n_1111),
	.B (n_831),
	.AN (n_813) );
   SEDFFX1 ar1_reg_13 ( .SI (ar1[12]),
	.SE (scan_en),
	.Q (ar1[13]),
	.E (n_4099),
	.D (\nbus_425[13] ),
	.CK (clk) );
   NAND3BX1 i_2254 ( .Y (n_1112),
	.C (n_869),
	.B (ir[0]),
	.AN (ir[2]) );
   SEDFFX1 ar1_reg_14 ( .SI (ar1[13]),
	.SE (scan_en),
	.Q (ar1[14]),
	.E (n_4099),
	.D (\nbus_425[14] ),
	.CK (clk) );
   SEDFFX1 ar1_reg_15 ( .SI (ar1[14]),
	.SE (scan_en),
	.Q (ar1[15]),
	.E (n_4099),
	.D (\nbus_425[15] ),
	.CK (clk) );
   NAND2BX1 i_2698 ( .Y (n_1114),
	.B (n_784),
	.AN (n_793) );
   INVX1 i_5175 ( .Y (n_4072),
	.A (n_1001) );
   INVX1 i_5176 ( .Y (n_4073),
	.A (n_998) );
   INVX1 i_5177 ( .Y (n_4074),
	.A (n_995) );
   INVX1 i_5178 ( .Y (n_4075),
	.A (n_1026) );
   INVX1 i_5179 ( .Y (n_4076),
	.A (n_922) );
   INVX1 i_5180 ( .Y (n_4077),
	.A (n_796) );
   INVX1 i_5181 ( .Y (n_4078),
	.A (n_820) );
   INVX1 i_5182 ( .Y (n_4079),
	.A (n_800) );
   INVX1 i_5183 ( .Y (n_4080),
	.A (n_801) );
   INVX1 i_5184 ( .Y (n_4081),
	.A (n_1111) );
   INVX1 i_5185 ( .Y (n_4082),
	.A (n_804) );
   INVX1 i_5186 ( .Y (n_4083),
	.A (n_1103) );
   INVX1 i_5187 ( .Y (n_4084),
	.A (n_790) );
   INVX1 i_5188 ( .Y (n_4085),
	.A (n_840) );
   INVX1 i_5189 ( .Y (n_4086),
	.A (n_872) );
   INVX1 i_5190 ( .Y (n_4087),
	.A (n_806) );
   INVX1 i_5191 ( .Y (n_4088),
	.A (n_816) );
   INVX1 i_5192 ( .Y (n_4089),
	.A (n_830) );
   INVX1 i_5193 ( .Y (n_4090),
	.A (n_784) );
   INVX1 i_5194 ( .Y (n_4091),
	.A (n_470) );
   INVX1 i_5195 ( .Y (n_4092),
	.A (two_cycle) );
   INVX1 i_5196 ( .Y (n_4093),
	.A (n_3128) );
   INVX1 i_5197 ( .Y (n_4094),
	.A (\nbus_440[0] ) );
   INVX1 i_5198 ( .Y (n_4095),
	.A (n_3742) );
   INVX1 i_5199 ( .Y (n_4096),
	.A (n_3748) );
   INVX1 i_5200 ( .Y (n_4097),
	.A (\nbus_428[0] ) );
   INVX1 i_5201 ( .Y (n_4098),
	.A (n_3976) );
   INVX1 i_5202 ( .Y (n_4099),
	.A (\nbus_424[0] ) );
   INVX1 i_5203 ( .Y (n_4100),
	.A (ir[8]) );
   INVX1 i_5204 ( .Y (n_4101),
	.A (pc[12]) );
   INVX1 i_5205 ( .Y (n_4220),
	.A (phi_1) );
   INVX1 i_5206 ( .Y (n_4221),
	.A (reset) );
   INVX1 i_5207 ( .Y (n_4222),
	.A (pc_acc) );
   INVX1 i_5208 ( .Y (n_4223),
	.A (ovm) );
   BUFX1 FE_OFC171_scan_enI ( .Y (FE_OFN171_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC166_scan_enI ( .Y (FE_OFN166_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC165_scan_enI ( .Y (FE_OFN165_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC164_scan_enI ( .Y (FE_OFN164_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC163_scan_enI ( .Y (FE_OFN163_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC162_scan_enI ( .Y (FE_OFN162_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC146_scan_enI ( .Y (FE_OFN146_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC145_scan_enI ( .Y (FE_OFN145_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC143_scan_enI ( .Y (FE_OFN143_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC142_scan_enI ( .Y (FE_OFN142_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC139_scan_enI ( .Y (FE_OFN139_scan_enI),
	.A (scan_en) );
   BUFX2 FE_OFC131_arp ( .Y (arp),
	.A (FE_OFN131_arp) );
   INVX2 FE_OFC130_dmov_inc ( .Y (dmov_inc),
	.A (FE_OFN130_dmov_inc) );
   INVXL FE_OFC129_dmov_inc ( .Y (FE_OFN130_dmov_inc),
	.A (FE_OFN129_dmov_inc) );
   BUFX1 FE_OFC17_scan_enI ( .Y (FE_OFN17_scan_enI),
	.A (FE_OFN145_scan_enI) );
   BUFX2 FE_OFC14_scan_enI ( .Y (FE_OFN14_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC13_scan_enI ( .Y (FE_OFN13_scan_enI),
	.A (scan_en) );
   BUFX2 FE_OFC9_scan_enI ( .Y (FE_OFN9_scan_enI),
	.A (FE_OFN139_scan_enI) );
endmodule

module m16x16 (
	a,
	b,
	y );
   input [15:0] a;
   input [15:0] b;
   output [31:0] y;

   // Internal wires
   wire n_465;
   wire n_447;
   wire n_1024;
   wire n_899;
   wire n_960;
   wire n_898;
   wire n_897;
   wire n_959;
   wire n_896;
   wire n_893;
   wire n_958;
   wire n_887;
   wire n_892;
   wire n_957;
   wire n_886;
   wire n_879;
   wire n_956;
   wire n_869;
   wire n_878;
   wire n_955;
   wire n_857;
   wire n_868;
   wire n_954;
   wire n_843;
   wire n_856;
   wire n_953;
   wire n_842;
   wire n_827;
   wire n_952;
   wire n_809;
   wire n_826;
   wire n_951;
   wire n_789;
   wire n_808;
   wire n_950;
   wire n_767;
   wire n_788;
   wire n_949;
   wire n_743;
   wire n_766;
   wire n_948;
   wire n_717;
   wire n_742;
   wire n_947;
   wire n_689;
   wire n_716;
   wire n_946;
   wire n_686;
   wire n_688;
   wire n_945;
   wire n_635;
   wire n_660;
   wire n_944;
   wire n_611;
   wire n_634;
   wire n_943;
   wire n_589;
   wire n_610;
   wire n_942;
   wire n_569;
   wire n_588;
   wire n_941;
   wire n_566;
   wire n_568;
   wire n_940;
   wire n_535;
   wire n_550;
   wire n_939;
   wire n_521;
   wire n_534;
   wire n_938;
   wire n_518;
   wire n_520;
   wire n_937;
   wire n_499;
   wire n_508;
   wire n_936;
   wire n_496;
   wire n_498;
   wire n_935;
   wire n_485;
   wire n_490;
   wire n_934;
   wire n_482;
   wire n_484;
   wire n_933;
   wire n_480;
   wire n_932;
   wire n_929;
   wire n_928;
   wire n_927;
   wire n_926;
   wire n_925;
   wire n_924;
   wire n_923;
   wire n_922;
   wire n_921;
   wire n_920;
   wire n_919;
   wire n_918;
   wire n_917;
   wire n_916;
   wire n_915;
   wire n_914;
   wire n_913;
   wire n_912;
   wire n_911;
   wire n_910;
   wire n_909;
   wire n_908;
   wire n_907;
   wire n_906;
   wire n_905;
   wire n_904;
   wire n_903;
   wire n_902;
   wire n_901;
   wire n_479;
   wire n_478;
   wire n_477;
   wire n_476;
   wire n_475;
   wire n_474;
   wire n_473;
   wire n_472;
   wire n_471;
   wire n_470;
   wire n_469;
   wire n_468;
   wire n_467;
   wire n_466;
   wire n_965;
   wire n_462;
   wire n_461;
   wire n_460;
   wire n_459;
   wire n_458;
   wire n_457;
   wire n_456;
   wire n_455;
   wire n_454;
   wire n_453;
   wire n_452;
   wire n_451;
   wire n_450;
   wire n_449;
   wire n_448;
   wire n_967;
   wire n_445;
   wire n_444;
   wire n_443;
   wire n_442;
   wire n_441;
   wire n_440;
   wire n_439;
   wire n_438;
   wire n_437;
   wire n_436;
   wire n_435;
   wire n_434;
   wire n_433;
   wire n_432;
   wire n_431;
   wire n_969;
   wire n_428;
   wire n_427;
   wire n_426;
   wire n_425;
   wire n_424;
   wire n_423;
   wire n_422;
   wire n_421;
   wire n_420;
   wire n_419;
   wire n_418;
   wire n_417;
   wire n_416;
   wire n_415;
   wire n_414;
   wire n_413;
   wire n_971;
   wire n_411;
   wire n_410;
   wire n_409;
   wire n_408;
   wire n_407;
   wire n_406;
   wire n_405;
   wire n_404;
   wire n_403;
   wire n_402;
   wire n_401;
   wire n_400;
   wire n_399;
   wire n_398;
   wire n_397;
   wire n_396;
   wire n_973;
   wire n_394;
   wire n_393;
   wire n_392;
   wire n_391;
   wire n_390;
   wire n_389;
   wire n_388;
   wire n_387;
   wire n_386;
   wire n_385;
   wire n_384;
   wire n_383;
   wire n_382;
   wire n_381;
   wire n_380;
   wire n_379;
   wire n_975;
   wire n_377;
   wire n_376;
   wire n_375;
   wire n_374;
   wire n_373;
   wire n_372;
   wire n_371;
   wire n_370;
   wire n_369;
   wire n_368;
   wire n_367;
   wire n_366;
   wire n_365;
   wire n_364;
   wire n_363;
   wire n_362;
   wire n_977;
   wire n_360;
   wire n_359;
   wire n_358;
   wire n_357;
   wire n_356;
   wire n_355;
   wire n_354;
   wire n_353;
   wire n_352;
   wire n_351;
   wire n_350;
   wire n_349;
   wire n_348;
   wire n_347;
   wire n_346;
   wire n_345;
   wire n_979;
   wire n_343;
   wire n_342;
   wire n_341;
   wire n_340;
   wire n_339;
   wire n_338;
   wire n_337;
   wire n_336;
   wire n_335;
   wire n_334;
   wire n_333;
   wire n_332;
   wire n_331;
   wire n_330;
   wire n_329;
   wire n_328;
   wire n_981;
   wire n_326;
   wire n_325;
   wire n_324;
   wire n_323;
   wire n_322;
   wire n_321;
   wire n_320;
   wire n_319;
   wire n_318;
   wire n_317;
   wire n_316;
   wire n_315;
   wire n_314;
   wire n_313;
   wire n_312;
   wire n_311;
   wire n_983;
   wire n_309;
   wire n_308;
   wire n_307;
   wire n_306;
   wire n_305;
   wire n_304;
   wire n_303;
   wire n_302;
   wire n_301;
   wire n_300;
   wire n_299;
   wire n_298;
   wire n_297;
   wire n_296;
   wire n_295;
   wire n_294;
   wire n_985;
   wire n_292;
   wire n_291;
   wire n_290;
   wire n_289;
   wire n_288;
   wire n_287;
   wire n_286;
   wire n_285;
   wire n_284;
   wire n_283;
   wire n_282;
   wire n_281;
   wire n_280;
   wire n_279;
   wire n_278;
   wire n_277;
   wire n_987;
   wire n_275;
   wire n_274;
   wire n_273;
   wire n_272;
   wire n_271;
   wire n_270;
   wire n_269;
   wire n_268;
   wire n_267;
   wire n_266;
   wire n_265;
   wire n_264;
   wire n_263;
   wire n_262;
   wire n_261;
   wire n_260;
   wire n_989;
   wire n_258;
   wire n_257;
   wire n_256;
   wire n_255;
   wire n_254;
   wire n_253;
   wire n_252;
   wire n_251;
   wire n_250;
   wire n_249;
   wire n_248;
   wire n_247;
   wire n_246;
   wire n_245;
   wire n_244;
   wire n_243;
   wire n_991;
   wire n_241;
   wire n_240;
   wire n_239;
   wire n_238;
   wire n_237;
   wire n_236;
   wire n_235;
   wire n_234;
   wire n_233;
   wire n_232;
   wire n_231;
   wire n_230;
   wire n_229;
   wire n_228;
   wire n_227;
   wire n_226;
   wire n_993;
   wire n_223;
   wire n_222;
   wire n_221;
   wire n_220;
   wire n_219;
   wire n_218;
   wire n_217;
   wire n_216;
   wire n_215;
   wire n_214;
   wire n_213;
   wire n_212;
   wire n_211;
   wire n_210;
   wire n_209;
   wire n_995;
   wire n_997;
   wire n_999;
   wire n_1001;
   wire n_1003;
   wire n_1005;
   wire n_1007;
   wire n_1009;
   wire n_1011;
   wire n_1013;
   wire n_1015;
   wire n_1017;
   wire n_1019;
   wire n_1021;
   wire n_1056;
   wire n_1057;
   wire n_1058;
   wire n_931;
   wire n_1059;
   wire n_1060;
   wire n_1061;
   wire n_1025;
   wire n_5393;
   wire n_1062;
   wire n_1063;
   wire n_1064;
   wire n_1086;
   wire n_1065;
   wire n_1066;
   wire n_1067;
   wire n_1087;
   wire n_1068;
   wire n_1069;
   wire n_1070;
   wire n_1148;
   wire n_5408;
   wire n_1071;
   wire n_1072;
   wire n_1073;
   wire n_1149;
   wire n_5413;
   wire n_1074;
   wire n_1075;
   wire n_1076;
   wire n_1150;
   wire n_5418;
   wire n_1077;
   wire n_1078;
   wire n_1079;
   wire n_1151;
   wire n_5423;
   wire n_1080;
   wire n_1081;
   wire n_1082;
   wire n_1212;
   wire n_1083;
   wire n_1118;
   wire n_1119;
   wire n_1213;
   wire n_1120;
   wire n_1121;
   wire n_1122;
   wire n_1214;
   wire n_1123;
   wire n_1124;
   wire n_1125;
   wire n_1215;
   wire n_1126;
   wire n_1127;
   wire n_1128;
   wire n_1216;
   wire n_1129;
   wire n_1130;
   wire n_1131;
   wire n_1217;
   wire n_1132;
   wire n_1133;
   wire n_1134;
   wire n_1218;
   wire n_1135;
   wire n_1136;
   wire n_1137;
   wire n_1219;
   wire n_1138;
   wire n_1139;
   wire n_1140;
   wire n_1280;
   wire n_5468;
   wire n_1141;
   wire n_1142;
   wire n_1143;
   wire n_1281;
   wire n_5473;
   wire n_1182;
   wire n_1183;
   wire n_1184;
   wire n_1282;
   wire n_5478;
   wire n_1185;
   wire n_1186;
   wire n_1187;
   wire n_1283;
   wire n_5483;
   wire n_1188;
   wire n_1189;
   wire n_1190;
   wire n_1284;
   wire n_5488;
   wire n_1191;
   wire n_1192;
   wire n_1193;
   wire n_1285;
   wire n_5493;
   wire n_1194;
   wire n_1195;
   wire n_1196;
   wire n_1286;
   wire n_5498;
   wire n_1197;
   wire n_1198;
   wire n_1199;
   wire n_1287;
   wire n_5503;
   wire n_1200;
   wire n_1201;
   wire n_1202;
   wire n_1288;
   wire n_5508;
   wire n_1203;
   wire n_1250;
   wire n_1251;
   wire n_1289;
   wire n_5513;
   wire n_1252;
   wire n_1253;
   wire n_1254;
   wire n_1290;
   wire n_5518;
   wire n_1255;
   wire n_1256;
   wire n_1257;
   wire n_1291;
   wire n_5523;
   wire n_1258;
   wire n_1259;
   wire n_1260;
   wire n_1292;
   wire n_5528;
   wire n_1261;
   wire n_1262;
   wire n_1263;
   wire n_1211;
   wire n_1210;
   wire n_1209;
   wire n_1208;
   wire n_1085;
   wire n_1147;
   wire n_1146;
   wire n_481;
   wire n_483;
   wire n_486;
   wire n_487;
   wire n_488;
   wire n_489;
   wire n_491;
   wire n_492;
   wire n_493;
   wire n_494;
   wire n_495;
   wire n_497;
   wire n_500;
   wire n_501;
   wire n_502;
   wire n_503;
   wire n_504;
   wire n_505;
   wire n_506;
   wire n_507;
   wire n_509;
   wire n_510;
   wire n_511;
   wire n_512;
   wire n_513;
   wire n_514;
   wire n_515;
   wire n_516;
   wire n_517;
   wire n_519;
   wire n_522;
   wire n_523;
   wire n_524;
   wire n_525;
   wire n_526;
   wire n_527;
   wire n_528;
   wire n_529;
   wire n_530;
   wire n_531;
   wire n_532;
   wire n_533;
   wire n_536;
   wire n_537;
   wire n_538;
   wire n_539;
   wire n_540;
   wire n_541;
   wire n_542;
   wire n_543;
   wire n_544;
   wire n_545;
   wire n_546;
   wire n_547;
   wire n_548;
   wire n_549;
   wire n_551;
   wire n_552;
   wire n_553;
   wire n_554;
   wire n_555;
   wire n_556;
   wire n_557;
   wire n_558;
   wire n_559;
   wire n_560;
   wire n_561;
   wire n_562;
   wire n_563;
   wire n_564;
   wire n_565;
   wire n_567;
   wire n_570;
   wire n_571;
   wire n_572;
   wire n_573;
   wire n_574;
   wire n_575;
   wire n_576;
   wire n_577;
   wire n_578;
   wire n_579;
   wire n_580;
   wire n_581;
   wire n_582;
   wire n_583;
   wire n_584;
   wire n_585;
   wire n_586;
   wire n_587;
   wire n_590;
   wire n_591;
   wire n_592;
   wire n_593;
   wire n_594;
   wire n_595;
   wire n_596;
   wire n_597;
   wire n_598;
   wire n_599;
   wire n_600;
   wire n_601;
   wire n_602;
   wire n_603;
   wire n_604;
   wire n_605;
   wire n_606;
   wire n_607;
   wire n_608;
   wire n_609;
   wire n_612;
   wire n_613;
   wire n_614;
   wire n_615;
   wire n_616;
   wire n_617;
   wire n_618;
   wire n_619;
   wire n_620;
   wire n_621;
   wire n_622;
   wire n_623;
   wire n_624;
   wire n_625;
   wire n_626;
   wire n_627;
   wire n_628;
   wire n_629;
   wire n_630;
   wire n_631;
   wire n_632;
   wire n_633;
   wire n_636;
   wire n_637;
   wire n_638;
   wire n_639;
   wire n_640;
   wire n_641;
   wire n_642;
   wire n_643;
   wire n_644;
   wire n_645;
   wire n_646;
   wire n_647;
   wire n_648;
   wire n_649;
   wire n_650;
   wire n_651;
   wire n_652;
   wire n_653;
   wire n_654;
   wire n_655;
   wire n_656;
   wire n_657;
   wire n_658;
   wire n_659;
   wire n_661;
   wire n_662;
   wire n_663;
   wire n_664;
   wire n_665;
   wire n_666;
   wire n_667;
   wire n_668;
   wire n_669;
   wire n_670;
   wire n_671;
   wire n_672;
   wire n_673;
   wire n_674;
   wire n_675;
   wire n_676;
   wire n_677;
   wire n_678;
   wire n_679;
   wire n_680;
   wire n_681;
   wire n_682;
   wire n_683;
   wire n_684;
   wire n_685;
   wire n_687;
   wire n_690;
   wire n_691;
   wire n_692;
   wire n_693;
   wire n_694;
   wire n_695;
   wire n_696;
   wire n_697;
   wire n_698;
   wire n_699;
   wire n_700;
   wire n_701;
   wire n_702;
   wire n_703;
   wire n_704;
   wire n_705;
   wire n_706;
   wire n_707;
   wire n_708;
   wire n_709;
   wire n_710;
   wire n_711;
   wire n_712;
   wire n_713;
   wire n_714;
   wire n_715;
   wire n_718;
   wire n_719;
   wire n_720;
   wire n_721;
   wire n_722;
   wire n_723;
   wire n_724;
   wire n_725;
   wire n_726;
   wire n_727;
   wire n_728;
   wire n_729;
   wire n_730;
   wire n_731;
   wire n_732;
   wire n_733;
   wire n_734;
   wire n_735;
   wire n_736;
   wire n_737;
   wire n_738;
   wire n_739;
   wire n_740;
   wire n_741;
   wire n_744;
   wire n_745;
   wire n_746;
   wire n_747;
   wire n_748;
   wire n_749;
   wire n_750;
   wire n_751;
   wire n_752;
   wire n_753;
   wire n_754;
   wire n_755;
   wire n_756;
   wire n_757;
   wire n_758;
   wire n_759;
   wire n_760;
   wire n_761;
   wire n_762;
   wire n_763;
   wire n_764;
   wire n_765;
   wire n_768;
   wire n_769;
   wire n_770;
   wire n_771;
   wire n_772;
   wire n_773;
   wire n_774;
   wire n_775;
   wire n_776;
   wire n_777;
   wire n_778;
   wire n_779;
   wire n_780;
   wire n_781;
   wire n_782;
   wire n_783;
   wire n_784;
   wire n_785;
   wire n_786;
   wire n_787;
   wire n_790;
   wire n_791;
   wire n_792;
   wire n_793;
   wire n_794;
   wire n_795;
   wire n_796;
   wire n_797;
   wire n_798;
   wire n_799;
   wire n_800;
   wire n_801;
   wire n_802;
   wire n_803;
   wire n_804;
   wire n_805;
   wire n_806;
   wire n_807;
   wire n_810;
   wire n_811;
   wire n_812;
   wire n_813;
   wire n_814;
   wire n_815;
   wire n_816;
   wire n_817;
   wire n_818;
   wire n_819;
   wire n_820;
   wire n_821;
   wire n_822;
   wire n_823;
   wire n_824;
   wire n_825;
   wire n_828;
   wire n_829;
   wire n_830;
   wire n_831;
   wire n_832;
   wire n_833;
   wire n_834;
   wire n_835;
   wire n_836;
   wire n_837;
   wire n_838;
   wire n_839;
   wire n_840;
   wire n_841;
   wire n_844;
   wire n_845;
   wire n_846;
   wire n_847;
   wire n_848;
   wire n_849;
   wire n_850;
   wire n_851;
   wire n_852;
   wire n_853;
   wire n_854;
   wire n_855;
   wire n_858;
   wire n_859;
   wire n_860;
   wire n_861;
   wire n_862;
   wire n_863;
   wire n_864;
   wire n_865;
   wire n_866;
   wire n_867;
   wire n_870;
   wire n_871;
   wire n_872;
   wire n_873;
   wire n_874;
   wire n_875;
   wire n_876;
   wire n_877;
   wire n_880;
   wire n_881;
   wire n_882;
   wire n_883;
   wire n_884;
   wire n_885;
   wire n_888;
   wire n_889;
   wire n_890;
   wire n_891;
   wire n_894;
   wire n_895;
   wire n_1026;
   wire n_1027;
   wire n_1028;
   wire n_1029;
   wire n_1030;
   wire n_1031;
   wire n_1032;
   wire n_1033;
   wire n_1034;
   wire n_1035;
   wire n_1036;
   wire n_1037;
   wire n_1038;
   wire n_1039;
   wire n_1040;
   wire n_1041;
   wire n_1042;
   wire n_1043;
   wire n_1044;
   wire n_1045;
   wire n_1046;
   wire n_1047;
   wire n_1048;
   wire n_1049;
   wire n_1050;
   wire n_1051;
   wire n_1052;
   wire n_1053;
   wire n_1088;
   wire n_1089;
   wire n_1090;
   wire n_1091;
   wire n_1092;
   wire n_1093;
   wire n_1094;
   wire n_1095;
   wire n_1096;
   wire n_1097;
   wire n_1098;
   wire n_1099;
   wire n_1100;
   wire n_1101;
   wire n_1102;
   wire n_1103;
   wire n_1104;
   wire n_1105;
   wire n_1106;
   wire n_1107;
   wire n_1108;
   wire n_1109;
   wire n_1110;
   wire n_1111;
   wire n_1112;
   wire n_1113;
   wire n_1152;
   wire n_1153;
   wire n_1154;
   wire n_1155;
   wire n_1156;
   wire n_1157;
   wire n_1158;
   wire n_1159;
   wire n_1160;
   wire n_1161;
   wire n_1162;
   wire n_1163;
   wire n_1164;
   wire n_1165;
   wire n_1166;
   wire n_1167;
   wire n_1168;
   wire n_1169;
   wire n_1170;
   wire n_1171;
   wire n_1172;
   wire n_1173;
   wire n_1220;
   wire n_1221;
   wire n_1222;
   wire n_1223;
   wire n_1224;
   wire n_1225;
   wire n_1226;
   wire n_1227;
   wire n_1228;
   wire n_1229;
   wire n_1230;
   wire n_1231;
   wire n_1232;
   wire n_1233;

   AOI21X1 i_561 ( .Y (y[1]),
	.B0 (n_1024),
	.A1 (n_447),
	.A0 (n_465) );
   NAND3X1 i_558 ( .Y (n_960),
	.C (n_899),
	.B (a[15]),
	.A (b[15]) );
   NAND2X1 i_557 ( .Y (n_959),
	.B (n_897),
	.A (n_898) );
   NAND2X1 i_556 ( .Y (n_958),
	.B (n_893),
	.A (n_896) );
   NAND2X1 i_555 ( .Y (n_957),
	.B (n_892),
	.A (n_887) );
   NAND2X1 i_554 ( .Y (n_956),
	.B (n_879),
	.A (n_886) );
   NAND2X1 i_553 ( .Y (n_955),
	.B (n_878),
	.A (n_869) );
   NAND2X1 i_552 ( .Y (n_954),
	.B (n_868),
	.A (n_857) );
   NAND2X1 i_551 ( .Y (n_953),
	.B (n_856),
	.A (n_843) );
   NAND2X1 i_550 ( .Y (n_952),
	.B (n_827),
	.A (n_842) );
   NAND2X1 i_549 ( .Y (n_951),
	.B (n_826),
	.A (n_809) );
   NAND2X1 i_548 ( .Y (n_950),
	.B (n_808),
	.A (n_789) );
   NAND2X1 i_547 ( .Y (n_949),
	.B (n_788),
	.A (n_767) );
   NAND2X1 i_546 ( .Y (n_948),
	.B (n_766),
	.A (n_743) );
   NAND2X1 i_545 ( .Y (n_947),
	.B (n_742),
	.A (n_717) );
   NAND2X1 i_544 ( .Y (n_946),
	.B (n_716),
	.A (n_689) );
   NAND2X1 i_543 ( .Y (n_945),
	.B (n_688),
	.A (n_686) );
   NAND2X1 i_542 ( .Y (n_944),
	.B (n_660),
	.A (n_635) );
   NAND2X1 i_541 ( .Y (n_943),
	.B (n_634),
	.A (n_611) );
   NAND2X1 i_540 ( .Y (n_942),
	.B (n_610),
	.A (n_589) );
   NAND2X1 i_539 ( .Y (n_941),
	.B (n_588),
	.A (n_569) );
   NAND2X1 i_538 ( .Y (n_940),
	.B (n_568),
	.A (n_566) );
   NAND2X1 i_537 ( .Y (n_939),
	.B (n_550),
	.A (n_535) );
   NAND2X1 i_536 ( .Y (n_938),
	.B (n_534),
	.A (n_521) );
   NAND2X1 i_535 ( .Y (n_937),
	.B (n_520),
	.A (n_518) );
   NAND2X1 i_534 ( .Y (n_936),
	.B (n_508),
	.A (n_499) );
   NAND2X1 i_533 ( .Y (n_935),
	.B (n_498),
	.A (n_496) );
   NAND2X1 i_532 ( .Y (n_934),
	.B (n_490),
	.A (n_485) );
   NAND2X1 i_531 ( .Y (n_933),
	.B (n_484),
	.A (n_482) );
   NAND3X1 i_530 ( .Y (n_932),
	.C (n_480),
	.B (a[0]),
	.A (b[2]) );
   NOR2X1 i_529 ( .Y (n_1024),
	.B (n_447),
	.A (n_465) );
   AOI21X1 i_527 ( .Y (n_929),
	.B0 (n_899),
	.A1 (a[15]),
	.A0 (b[15]) );
   NOR2X1 i_526 ( .Y (n_928),
	.B (n_897),
	.A (n_898) );
   NOR2X1 i_525 ( .Y (n_927),
	.B (n_893),
	.A (n_896) );
   NOR2X1 i_524 ( .Y (n_926),
	.B (n_892),
	.A (n_887) );
   NOR2X1 i_523 ( .Y (n_925),
	.B (n_879),
	.A (n_886) );
   NOR2X1 i_522 ( .Y (n_924),
	.B (n_878),
	.A (n_869) );
   NOR2X1 i_521 ( .Y (n_923),
	.B (n_868),
	.A (n_857) );
   NOR2X1 i_520 ( .Y (n_922),
	.B (n_856),
	.A (n_843) );
   NOR2X1 i_519 ( .Y (n_921),
	.B (n_827),
	.A (n_842) );
   NOR2X1 i_518 ( .Y (n_920),
	.B (n_826),
	.A (n_809) );
   NOR2X1 i_517 ( .Y (n_919),
	.B (n_808),
	.A (n_789) );
   NOR2X1 i_516 ( .Y (n_918),
	.B (n_788),
	.A (n_767) );
   NOR2X1 i_515 ( .Y (n_917),
	.B (n_766),
	.A (n_743) );
   NOR2X1 i_514 ( .Y (n_916),
	.B (n_742),
	.A (n_717) );
   NOR2X1 i_513 ( .Y (n_915),
	.B (n_716),
	.A (n_689) );
   NOR2X1 i_512 ( .Y (n_914),
	.B (n_688),
	.A (n_686) );
   NOR2X1 i_511 ( .Y (n_913),
	.B (n_660),
	.A (n_635) );
   NOR2X1 i_510 ( .Y (n_912),
	.B (n_634),
	.A (n_611) );
   NOR2X1 i_509 ( .Y (n_911),
	.B (n_610),
	.A (n_589) );
   NOR2X1 i_508 ( .Y (n_910),
	.B (n_588),
	.A (n_569) );
   NOR2X1 i_507 ( .Y (n_909),
	.B (n_568),
	.A (n_566) );
   NOR2X1 i_506 ( .Y (n_908),
	.B (n_550),
	.A (n_535) );
   NOR2X1 i_505 ( .Y (n_907),
	.B (n_534),
	.A (n_521) );
   NOR2X1 i_504 ( .Y (n_906),
	.B (n_520),
	.A (n_518) );
   NOR2X1 i_503 ( .Y (n_905),
	.B (n_508),
	.A (n_499) );
   NOR2X1 i_502 ( .Y (n_904),
	.B (n_498),
	.A (n_496) );
   NOR2X1 i_501 ( .Y (n_903),
	.B (n_490),
	.A (n_485) );
   NOR2X1 i_500 ( .Y (n_902),
	.B (n_484),
	.A (n_482) );
   AOI21X1 i_499 ( .Y (n_901),
	.B0 (n_480),
	.A1 (a[0]),
	.A0 (b[2]) );
   AND2X1 i_287 ( .Y (n_479),
	.B (a[15]),
	.A (b[0]) );
   AND2X1 i_286 ( .Y (n_478),
	.B (a[14]),
	.A (b[0]) );
   AND2X1 i_285 ( .Y (n_477),
	.B (a[13]),
	.A (b[0]) );
   AND2X1 i_284 ( .Y (n_476),
	.B (a[12]),
	.A (b[0]) );
   AND2X1 i_283 ( .Y (n_475),
	.B (a[11]),
	.A (b[0]) );
   AND2X1 i_282 ( .Y (n_474),
	.B (a[10]),
	.A (b[0]) );
   AND2X1 i_281 ( .Y (n_473),
	.B (a[9]),
	.A (b[0]) );
   AND2X1 i_280 ( .Y (n_472),
	.B (a[8]),
	.A (b[0]) );
   AND2X1 i_279 ( .Y (n_471),
	.B (a[7]),
	.A (b[0]) );
   AND2X1 i_278 ( .Y (n_470),
	.B (a[6]),
	.A (b[0]) );
   AND2X1 i_277 ( .Y (n_469),
	.B (a[5]),
	.A (b[0]) );
   AND2X1 i_276 ( .Y (n_468),
	.B (a[4]),
	.A (b[0]) );
   AND2X1 i_275 ( .Y (n_467),
	.B (a[3]),
	.A (b[0]) );
   AND2X1 i_274 ( .Y (n_466),
	.B (a[2]),
	.A (b[0]) );
   NAND2X1 i_273 ( .Y (n_465),
	.B (a[1]),
	.A (b[0]) );
   AND2X1 i_272 ( .Y (y[0]),
	.B (a[0]),
	.A (b[0]) );
   AOI31X1 i_563 ( .Y (n_965),
	.B0 (n_901),
	.A2 (n_480),
	.A1 (a[0]),
	.A0 (b[2]) );
   AND2X1 i_270 ( .Y (n_462),
	.B (a[15]),
	.A (b[1]) );
   AND2X1 i_269 ( .Y (n_461),
	.B (a[14]),
	.A (b[1]) );
   AND2X1 i_268 ( .Y (n_460),
	.B (a[13]),
	.A (b[1]) );
   AND2X1 i_267 ( .Y (n_459),
	.B (a[12]),
	.A (b[1]) );
   AND2X1 i_266 ( .Y (n_458),
	.B (a[11]),
	.A (b[1]) );
   AND2X1 i_265 ( .Y (n_457),
	.B (a[10]),
	.A (b[1]) );
   AND2X1 i_264 ( .Y (n_456),
	.B (a[9]),
	.A (b[1]) );
   AND2X1 i_263 ( .Y (n_455),
	.B (a[8]),
	.A (b[1]) );
   AND2X1 i_262 ( .Y (n_454),
	.B (a[7]),
	.A (b[1]) );
   AND2X1 i_261 ( .Y (n_453),
	.B (a[6]),
	.A (b[1]) );
   AND2X1 i_260 ( .Y (n_452),
	.B (a[5]),
	.A (b[1]) );
   AND2X1 i_259 ( .Y (n_451),
	.B (a[4]),
	.A (b[1]) );
   AND2X1 i_258 ( .Y (n_450),
	.B (a[3]),
	.A (b[1]) );
   AND2X1 i_257 ( .Y (n_449),
	.B (a[2]),
	.A (b[1]) );
   AND2X1 i_256 ( .Y (n_448),
	.B (a[1]),
	.A (b[1]) );
   NAND2X1 i_255 ( .Y (n_447),
	.B (a[0]),
	.A (b[1]) );
   AOI21X1 i_565 ( .Y (n_967),
	.B0 (n_902),
	.A1 (n_484),
	.A0 (n_482) );
   AND2X1 i_253 ( .Y (n_445),
	.B (a[15]),
	.A (b[2]) );
   AND2X1 i_252 ( .Y (n_444),
	.B (a[14]),
	.A (b[2]) );
   AND2X1 i_251 ( .Y (n_443),
	.B (a[13]),
	.A (b[2]) );
   AND2X1 i_250 ( .Y (n_442),
	.B (a[12]),
	.A (b[2]) );
   AND2X1 i_249 ( .Y (n_441),
	.B (a[11]),
	.A (b[2]) );
   AND2X1 i_248 ( .Y (n_440),
	.B (a[10]),
	.A (b[2]) );
   AND2X1 i_247 ( .Y (n_439),
	.B (a[9]),
	.A (b[2]) );
   AND2X1 i_246 ( .Y (n_438),
	.B (a[8]),
	.A (b[2]) );
   AND2X1 i_245 ( .Y (n_437),
	.B (a[7]),
	.A (b[2]) );
   AND2X1 i_244 ( .Y (n_436),
	.B (a[6]),
	.A (b[2]) );
   AND2X1 i_243 ( .Y (n_435),
	.B (a[5]),
	.A (b[2]) );
   AND2X1 i_242 ( .Y (n_434),
	.B (a[4]),
	.A (b[2]) );
   AND2X1 i_241 ( .Y (n_433),
	.B (a[3]),
	.A (b[2]) );
   AND2X1 i_240 ( .Y (n_432),
	.B (a[2]),
	.A (b[2]) );
   AND2X1 i_239 ( .Y (n_431),
	.B (a[1]),
	.A (b[2]) );
   AOI21X1 i_567 ( .Y (n_969),
	.B0 (n_903),
	.A1 (n_490),
	.A0 (n_485) );
   AND2X1 i_236 ( .Y (n_428),
	.B (a[15]),
	.A (b[3]) );
   AND2X1 i_235 ( .Y (n_427),
	.B (a[14]),
	.A (b[3]) );
   AND2X1 i_234 ( .Y (n_426),
	.B (a[13]),
	.A (b[3]) );
   AND2X1 i_233 ( .Y (n_425),
	.B (a[12]),
	.A (b[3]) );
   AND2X1 i_232 ( .Y (n_424),
	.B (a[11]),
	.A (b[3]) );
   AND2X1 i_231 ( .Y (n_423),
	.B (a[10]),
	.A (b[3]) );
   AND2X1 i_230 ( .Y (n_422),
	.B (a[9]),
	.A (b[3]) );
   AND2X1 i_229 ( .Y (n_421),
	.B (a[8]),
	.A (b[3]) );
   AND2X1 i_228 ( .Y (n_420),
	.B (a[7]),
	.A (b[3]) );
   AND2X1 i_227 ( .Y (n_419),
	.B (a[6]),
	.A (b[3]) );
   AND2X1 i_226 ( .Y (n_418),
	.B (a[5]),
	.A (b[3]) );
   AND2X1 i_225 ( .Y (n_417),
	.B (a[4]),
	.A (b[3]) );
   AND2X1 i_224 ( .Y (n_416),
	.B (a[3]),
	.A (b[3]) );
   AND2X1 i_223 ( .Y (n_415),
	.B (a[2]),
	.A (b[3]) );
   AND2X1 i_222 ( .Y (n_414),
	.B (a[1]),
	.A (b[3]) );
   AND2X1 i_221 ( .Y (n_413),
	.B (a[0]),
	.A (b[3]) );
   AOI21X1 i_569 ( .Y (n_971),
	.B0 (n_904),
	.A1 (n_498),
	.A0 (n_496) );
   AND2X1 i_219 ( .Y (n_411),
	.B (a[15]),
	.A (b[4]) );
   AND2X1 i_218 ( .Y (n_410),
	.B (a[14]),
	.A (b[4]) );
   AND2X1 i_217 ( .Y (n_409),
	.B (a[13]),
	.A (b[4]) );
   AND2X1 i_216 ( .Y (n_408),
	.B (a[12]),
	.A (b[4]) );
   AND2X1 i_215 ( .Y (n_407),
	.B (a[11]),
	.A (b[4]) );
   AND2X1 i_214 ( .Y (n_406),
	.B (a[10]),
	.A (b[4]) );
   AND2X1 i_213 ( .Y (n_405),
	.B (a[9]),
	.A (b[4]) );
   AND2X1 i_212 ( .Y (n_404),
	.B (a[8]),
	.A (b[4]) );
   AND2X1 i_211 ( .Y (n_403),
	.B (a[7]),
	.A (b[4]) );
   AND2X1 i_210 ( .Y (n_402),
	.B (a[6]),
	.A (b[4]) );
   AND2X1 i_209 ( .Y (n_401),
	.B (a[5]),
	.A (b[4]) );
   AND2X1 i_208 ( .Y (n_400),
	.B (a[4]),
	.A (b[4]) );
   AND2X1 i_207 ( .Y (n_399),
	.B (a[3]),
	.A (b[4]) );
   AND2X1 i_206 ( .Y (n_398),
	.B (a[2]),
	.A (b[4]) );
   AND2X1 i_205 ( .Y (n_397),
	.B (a[1]),
	.A (b[4]) );
   AND2X1 i_204 ( .Y (n_396),
	.B (a[0]),
	.A (b[4]) );
   AOI21X1 i_571 ( .Y (n_973),
	.B0 (n_905),
	.A1 (n_508),
	.A0 (n_499) );
   AND2X1 i_202 ( .Y (n_394),
	.B (a[15]),
	.A (b[5]) );
   AND2X1 i_201 ( .Y (n_393),
	.B (a[14]),
	.A (b[5]) );
   AND2X1 i_200 ( .Y (n_392),
	.B (a[13]),
	.A (b[5]) );
   AND2X1 i_199 ( .Y (n_391),
	.B (a[12]),
	.A (b[5]) );
   AND2X1 i_198 ( .Y (n_390),
	.B (a[11]),
	.A (b[5]) );
   AND2X1 i_197 ( .Y (n_389),
	.B (a[10]),
	.A (b[5]) );
   AND2X1 i_196 ( .Y (n_388),
	.B (a[9]),
	.A (b[5]) );
   AND2X1 i_195 ( .Y (n_387),
	.B (a[8]),
	.A (b[5]) );
   AND2X1 i_194 ( .Y (n_386),
	.B (a[7]),
	.A (b[5]) );
   AND2X1 i_193 ( .Y (n_385),
	.B (a[6]),
	.A (b[5]) );
   AND2X1 i_192 ( .Y (n_384),
	.B (a[5]),
	.A (b[5]) );
   AND2X1 i_191 ( .Y (n_383),
	.B (a[4]),
	.A (b[5]) );
   AND2X1 i_190 ( .Y (n_382),
	.B (a[3]),
	.A (b[5]) );
   AND2X1 i_189 ( .Y (n_381),
	.B (a[2]),
	.A (b[5]) );
   AND2X1 i_188 ( .Y (n_380),
	.B (a[1]),
	.A (b[5]) );
   AND2X1 i_187 ( .Y (n_379),
	.B (a[0]),
	.A (b[5]) );
   AOI21X1 i_573 ( .Y (n_975),
	.B0 (n_906),
	.A1 (n_520),
	.A0 (n_518) );
   AND2X1 i_185 ( .Y (n_377),
	.B (a[15]),
	.A (b[6]) );
   AND2X1 i_184 ( .Y (n_376),
	.B (a[14]),
	.A (b[6]) );
   AND2X1 i_183 ( .Y (n_375),
	.B (a[13]),
	.A (b[6]) );
   AND2X1 i_182 ( .Y (n_374),
	.B (a[12]),
	.A (b[6]) );
   AND2X1 i_181 ( .Y (n_373),
	.B (a[11]),
	.A (b[6]) );
   AND2X1 i_180 ( .Y (n_372),
	.B (a[10]),
	.A (b[6]) );
   AND2X1 i_179 ( .Y (n_371),
	.B (a[9]),
	.A (b[6]) );
   AND2X1 i_178 ( .Y (n_370),
	.B (a[8]),
	.A (b[6]) );
   AND2X1 i_177 ( .Y (n_369),
	.B (a[7]),
	.A (b[6]) );
   AND2X1 i_176 ( .Y (n_368),
	.B (a[6]),
	.A (b[6]) );
   AND2X1 i_175 ( .Y (n_367),
	.B (a[5]),
	.A (b[6]) );
   AND2X1 i_174 ( .Y (n_366),
	.B (a[4]),
	.A (b[6]) );
   AND2X1 i_173 ( .Y (n_365),
	.B (a[3]),
	.A (b[6]) );
   AND2X1 i_172 ( .Y (n_364),
	.B (a[2]),
	.A (b[6]) );
   AND2X1 i_171 ( .Y (n_363),
	.B (a[1]),
	.A (b[6]) );
   AND2X1 i_170 ( .Y (n_362),
	.B (a[0]),
	.A (b[6]) );
   AOI21X1 i_575 ( .Y (n_977),
	.B0 (n_907),
	.A1 (n_534),
	.A0 (n_521) );
   AND2X1 i_168 ( .Y (n_360),
	.B (a[15]),
	.A (b[7]) );
   AND2X1 i_167 ( .Y (n_359),
	.B (a[14]),
	.A (b[7]) );
   AND2X1 i_166 ( .Y (n_358),
	.B (a[13]),
	.A (b[7]) );
   AND2X1 i_165 ( .Y (n_357),
	.B (a[12]),
	.A (b[7]) );
   AND2X1 i_164 ( .Y (n_356),
	.B (a[11]),
	.A (b[7]) );
   AND2X1 i_163 ( .Y (n_355),
	.B (a[10]),
	.A (b[7]) );
   AND2X1 i_162 ( .Y (n_354),
	.B (a[9]),
	.A (b[7]) );
   AND2X1 i_161 ( .Y (n_353),
	.B (a[8]),
	.A (b[7]) );
   AND2X1 i_160 ( .Y (n_352),
	.B (a[7]),
	.A (b[7]) );
   AND2X1 i_159 ( .Y (n_351),
	.B (a[6]),
	.A (b[7]) );
   AND2X1 i_158 ( .Y (n_350),
	.B (a[5]),
	.A (b[7]) );
   AND2X1 i_157 ( .Y (n_349),
	.B (a[4]),
	.A (b[7]) );
   AND2X1 i_156 ( .Y (n_348),
	.B (a[3]),
	.A (b[7]) );
   AND2X1 i_155 ( .Y (n_347),
	.B (a[2]),
	.A (b[7]) );
   AND2X1 i_154 ( .Y (n_346),
	.B (a[1]),
	.A (b[7]) );
   AND2X1 i_153 ( .Y (n_345),
	.B (a[0]),
	.A (b[7]) );
   AOI21X1 i_577 ( .Y (n_979),
	.B0 (n_908),
	.A1 (n_550),
	.A0 (n_535) );
   AND2X1 i_151 ( .Y (n_343),
	.B (a[15]),
	.A (b[8]) );
   AND2X1 i_150 ( .Y (n_342),
	.B (a[14]),
	.A (b[8]) );
   AND2X1 i_149 ( .Y (n_341),
	.B (a[13]),
	.A (b[8]) );
   AND2X1 i_148 ( .Y (n_340),
	.B (a[12]),
	.A (b[8]) );
   AND2X1 i_147 ( .Y (n_339),
	.B (a[11]),
	.A (b[8]) );
   AND2X1 i_146 ( .Y (n_338),
	.B (a[10]),
	.A (b[8]) );
   AND2X1 i_145 ( .Y (n_337),
	.B (a[9]),
	.A (b[8]) );
   AND2X1 i_144 ( .Y (n_336),
	.B (a[8]),
	.A (b[8]) );
   AND2X1 i_143 ( .Y (n_335),
	.B (a[7]),
	.A (b[8]) );
   AND2X1 i_142 ( .Y (n_334),
	.B (a[6]),
	.A (b[8]) );
   AND2X1 i_141 ( .Y (n_333),
	.B (a[5]),
	.A (b[8]) );
   AND2X1 i_140 ( .Y (n_332),
	.B (a[4]),
	.A (b[8]) );
   AND2X1 i_139 ( .Y (n_331),
	.B (a[3]),
	.A (b[8]) );
   AND2X1 i_138 ( .Y (n_330),
	.B (a[2]),
	.A (b[8]) );
   AND2X1 i_137 ( .Y (n_329),
	.B (a[1]),
	.A (b[8]) );
   AND2X1 i_136 ( .Y (n_328),
	.B (a[0]),
	.A (b[8]) );
   AOI21X1 i_579 ( .Y (n_981),
	.B0 (n_909),
	.A1 (n_568),
	.A0 (n_566) );
   AND2X1 i_134 ( .Y (n_326),
	.B (a[15]),
	.A (b[9]) );
   AND2X1 i_133 ( .Y (n_325),
	.B (a[14]),
	.A (b[9]) );
   AND2X1 i_132 ( .Y (n_324),
	.B (a[13]),
	.A (b[9]) );
   AND2X1 i_131 ( .Y (n_323),
	.B (a[12]),
	.A (b[9]) );
   AND2X1 i_130 ( .Y (n_322),
	.B (a[11]),
	.A (b[9]) );
   AND2X1 i_129 ( .Y (n_321),
	.B (a[10]),
	.A (b[9]) );
   AND2X1 i_128 ( .Y (n_320),
	.B (a[9]),
	.A (b[9]) );
   AND2X1 i_127 ( .Y (n_319),
	.B (a[8]),
	.A (b[9]) );
   AND2X1 i_126 ( .Y (n_318),
	.B (a[7]),
	.A (b[9]) );
   AND2X1 i_125 ( .Y (n_317),
	.B (a[6]),
	.A (b[9]) );
   AND2X1 i_124 ( .Y (n_316),
	.B (a[5]),
	.A (b[9]) );
   AND2X1 i_123 ( .Y (n_315),
	.B (a[4]),
	.A (b[9]) );
   AND2X1 i_122 ( .Y (n_314),
	.B (a[3]),
	.A (b[9]) );
   AND2X1 i_121 ( .Y (n_313),
	.B (a[2]),
	.A (b[9]) );
   AND2X1 i_120 ( .Y (n_312),
	.B (a[1]),
	.A (b[9]) );
   AND2X1 i_119 ( .Y (n_311),
	.B (a[0]),
	.A (b[9]) );
   AOI21X1 i_581 ( .Y (n_983),
	.B0 (n_910),
	.A1 (n_588),
	.A0 (n_569) );
   AND2X1 i_117 ( .Y (n_309),
	.B (a[15]),
	.A (b[10]) );
   AND2X1 i_116 ( .Y (n_308),
	.B (a[14]),
	.A (b[10]) );
   AND2X1 i_115 ( .Y (n_307),
	.B (a[13]),
	.A (b[10]) );
   AND2X1 i_114 ( .Y (n_306),
	.B (a[12]),
	.A (b[10]) );
   AND2X1 i_113 ( .Y (n_305),
	.B (a[11]),
	.A (b[10]) );
   AND2X1 i_112 ( .Y (n_304),
	.B (a[10]),
	.A (b[10]) );
   AND2X1 i_111 ( .Y (n_303),
	.B (a[9]),
	.A (b[10]) );
   AND2X1 i_110 ( .Y (n_302),
	.B (a[8]),
	.A (b[10]) );
   AND2X1 i_109 ( .Y (n_301),
	.B (a[7]),
	.A (b[10]) );
   AND2X1 i_108 ( .Y (n_300),
	.B (a[6]),
	.A (b[10]) );
   AND2X1 i_107 ( .Y (n_299),
	.B (a[5]),
	.A (b[10]) );
   AND2X1 i_106 ( .Y (n_298),
	.B (a[4]),
	.A (b[10]) );
   AND2X1 i_105 ( .Y (n_297),
	.B (a[3]),
	.A (b[10]) );
   AND2X1 i_104 ( .Y (n_296),
	.B (a[2]),
	.A (b[10]) );
   AND2X1 i_103 ( .Y (n_295),
	.B (a[1]),
	.A (b[10]) );
   AND2X1 i_102 ( .Y (n_294),
	.B (a[0]),
	.A (b[10]) );
   AOI21X1 i_583 ( .Y (n_985),
	.B0 (n_911),
	.A1 (n_610),
	.A0 (n_589) );
   AND2X1 i_100 ( .Y (n_292),
	.B (a[15]),
	.A (b[11]) );
   AND2X1 i_99 ( .Y (n_291),
	.B (a[14]),
	.A (b[11]) );
   AND2X1 i_98 ( .Y (n_290),
	.B (a[13]),
	.A (b[11]) );
   AND2X1 i_97 ( .Y (n_289),
	.B (a[12]),
	.A (b[11]) );
   AND2X1 i_96 ( .Y (n_288),
	.B (a[11]),
	.A (b[11]) );
   AND2X1 i_95 ( .Y (n_287),
	.B (a[10]),
	.A (b[11]) );
   AND2X1 i_94 ( .Y (n_286),
	.B (a[9]),
	.A (b[11]) );
   AND2X1 i_93 ( .Y (n_285),
	.B (a[8]),
	.A (b[11]) );
   AND2X1 i_92 ( .Y (n_284),
	.B (a[7]),
	.A (b[11]) );
   AND2X1 i_91 ( .Y (n_283),
	.B (a[6]),
	.A (b[11]) );
   AND2X1 i_90 ( .Y (n_282),
	.B (a[5]),
	.A (b[11]) );
   AND2X1 i_89 ( .Y (n_281),
	.B (a[4]),
	.A (b[11]) );
   AND2X1 i_88 ( .Y (n_280),
	.B (a[3]),
	.A (b[11]) );
   AND2X1 i_87 ( .Y (n_279),
	.B (a[2]),
	.A (b[11]) );
   AND2X1 i_86 ( .Y (n_278),
	.B (a[1]),
	.A (b[11]) );
   AND2X1 i_85 ( .Y (n_277),
	.B (a[0]),
	.A (b[11]) );
   AOI21X1 i_585 ( .Y (n_987),
	.B0 (n_912),
	.A1 (n_634),
	.A0 (n_611) );
   AND2X1 i_83 ( .Y (n_275),
	.B (a[15]),
	.A (b[12]) );
   AND2X1 i_82 ( .Y (n_274),
	.B (a[14]),
	.A (b[12]) );
   AND2X1 i_81 ( .Y (n_273),
	.B (a[13]),
	.A (b[12]) );
   AND2X1 i_80 ( .Y (n_272),
	.B (a[12]),
	.A (b[12]) );
   AND2X1 i_79 ( .Y (n_271),
	.B (a[11]),
	.A (b[12]) );
   AND2X1 i_78 ( .Y (n_270),
	.B (a[10]),
	.A (b[12]) );
   AND2X1 i_77 ( .Y (n_269),
	.B (a[9]),
	.A (b[12]) );
   AND2X1 i_76 ( .Y (n_268),
	.B (a[8]),
	.A (b[12]) );
   AND2X1 i_75 ( .Y (n_267),
	.B (a[7]),
	.A (b[12]) );
   AND2X1 i_74 ( .Y (n_266),
	.B (a[6]),
	.A (b[12]) );
   AND2X1 i_73 ( .Y (n_265),
	.B (a[5]),
	.A (b[12]) );
   AND2X1 i_72 ( .Y (n_264),
	.B (a[4]),
	.A (b[12]) );
   AND2X1 i_71 ( .Y (n_263),
	.B (a[3]),
	.A (b[12]) );
   AND2X1 i_70 ( .Y (n_262),
	.B (a[2]),
	.A (b[12]) );
   AND2X1 i_69 ( .Y (n_261),
	.B (a[1]),
	.A (b[12]) );
   AND2X1 i_68 ( .Y (n_260),
	.B (a[0]),
	.A (b[12]) );
   AOI21X1 i_587 ( .Y (n_989),
	.B0 (n_913),
	.A1 (n_660),
	.A0 (n_635) );
   AND2X1 i_66 ( .Y (n_258),
	.B (a[15]),
	.A (b[13]) );
   AND2X1 i_65 ( .Y (n_257),
	.B (a[14]),
	.A (b[13]) );
   AND2X1 i_64 ( .Y (n_256),
	.B (a[13]),
	.A (b[13]) );
   AND2X1 i_63 ( .Y (n_255),
	.B (a[12]),
	.A (b[13]) );
   AND2X1 i_62 ( .Y (n_254),
	.B (a[11]),
	.A (b[13]) );
   AND2X1 i_61 ( .Y (n_253),
	.B (a[10]),
	.A (b[13]) );
   AND2X1 i_60 ( .Y (n_252),
	.B (a[9]),
	.A (b[13]) );
   AND2X1 i_59 ( .Y (n_251),
	.B (a[8]),
	.A (b[13]) );
   AND2X1 i_58 ( .Y (n_250),
	.B (a[7]),
	.A (b[13]) );
   AND2X1 i_57 ( .Y (n_249),
	.B (a[6]),
	.A (b[13]) );
   AND2X1 i_56 ( .Y (n_248),
	.B (a[5]),
	.A (b[13]) );
   AND2X1 i_55 ( .Y (n_247),
	.B (a[4]),
	.A (b[13]) );
   AND2X1 i_54 ( .Y (n_246),
	.B (a[3]),
	.A (b[13]) );
   AND2X1 i_53 ( .Y (n_245),
	.B (a[2]),
	.A (b[13]) );
   AND2X1 i_52 ( .Y (n_244),
	.B (a[1]),
	.A (b[13]) );
   AND2X1 i_51 ( .Y (n_243),
	.B (a[0]),
	.A (b[13]) );
   AOI21X1 i_589 ( .Y (n_991),
	.B0 (n_914),
	.A1 (n_688),
	.A0 (n_686) );
   AND2X1 i_49 ( .Y (n_241),
	.B (a[15]),
	.A (b[14]) );
   AND2X1 i_48 ( .Y (n_240),
	.B (a[14]),
	.A (b[14]) );
   AND2X1 i_47 ( .Y (n_239),
	.B (a[13]),
	.A (b[14]) );
   AND2X1 i_46 ( .Y (n_238),
	.B (a[12]),
	.A (b[14]) );
   AND2X1 i_45 ( .Y (n_237),
	.B (a[11]),
	.A (b[14]) );
   AND2X1 i_44 ( .Y (n_236),
	.B (a[10]),
	.A (b[14]) );
   AND2X1 i_43 ( .Y (n_235),
	.B (a[9]),
	.A (b[14]) );
   AND2X1 i_42 ( .Y (n_234),
	.B (a[8]),
	.A (b[14]) );
   AND2X1 i_41 ( .Y (n_233),
	.B (a[7]),
	.A (b[14]) );
   AND2X1 i_40 ( .Y (n_232),
	.B (a[6]),
	.A (b[14]) );
   AND2X1 i_39 ( .Y (n_231),
	.B (a[5]),
	.A (b[14]) );
   AND2X1 i_38 ( .Y (n_230),
	.B (a[4]),
	.A (b[14]) );
   AND2X1 i_37 ( .Y (n_229),
	.B (a[3]),
	.A (b[14]) );
   AND2X1 i_36 ( .Y (n_228),
	.B (a[2]),
	.A (b[14]) );
   AND2X1 i_35 ( .Y (n_227),
	.B (a[1]),
	.A (b[14]) );
   AND2X1 i_34 ( .Y (n_226),
	.B (a[0]),
	.A (b[14]) );
   AOI21X1 i_591 ( .Y (n_993),
	.B0 (n_915),
	.A1 (n_716),
	.A0 (n_689) );
   AND2X1 i_31 ( .Y (n_223),
	.B (a[14]),
	.A (b[15]) );
   AND2X1 i_30 ( .Y (n_222),
	.B (a[13]),
	.A (b[15]) );
   AND2X1 i_29 ( .Y (n_221),
	.B (a[12]),
	.A (b[15]) );
   AND2X1 i_28 ( .Y (n_220),
	.B (a[11]),
	.A (b[15]) );
   AND2X1 i_27 ( .Y (n_219),
	.B (a[10]),
	.A (b[15]) );
   AND2X1 i_26 ( .Y (n_218),
	.B (a[9]),
	.A (b[15]) );
   AND2X1 i_25 ( .Y (n_217),
	.B (a[8]),
	.A (b[15]) );
   AND2X1 i_24 ( .Y (n_216),
	.B (a[7]),
	.A (b[15]) );
   AND2X1 i_23 ( .Y (n_215),
	.B (a[6]),
	.A (b[15]) );
   AND2X1 i_22 ( .Y (n_214),
	.B (a[5]),
	.A (b[15]) );
   AND2X1 i_21 ( .Y (n_213),
	.B (a[4]),
	.A (b[15]) );
   AND2X1 i_20 ( .Y (n_212),
	.B (a[3]),
	.A (b[15]) );
   AND2X1 i_19 ( .Y (n_211),
	.B (a[2]),
	.A (b[15]) );
   AND2X1 i_18 ( .Y (n_210),
	.B (a[1]),
	.A (b[15]) );
   AND2X1 i_17 ( .Y (n_209),
	.B (a[0]),
	.A (b[15]) );
   AOI21X1 i_593 ( .Y (n_995),
	.B0 (n_916),
	.A1 (n_742),
	.A0 (n_717) );
   AOI21X1 i_595 ( .Y (n_997),
	.B0 (n_917),
	.A1 (n_766),
	.A0 (n_743) );
   AOI21X1 i_597 ( .Y (n_999),
	.B0 (n_918),
	.A1 (n_788),
	.A0 (n_767) );
   AOI21X1 i_599 ( .Y (n_1001),
	.B0 (n_919),
	.A1 (n_808),
	.A0 (n_789) );
   AOI21X1 i_601 ( .Y (n_1003),
	.B0 (n_920),
	.A1 (n_826),
	.A0 (n_809) );
   AOI21X1 i_603 ( .Y (n_1005),
	.B0 (n_921),
	.A1 (n_827),
	.A0 (n_842) );
   AOI21X1 i_605 ( .Y (n_1007),
	.B0 (n_922),
	.A1 (n_856),
	.A0 (n_843) );
   AOI21X1 i_607 ( .Y (n_1009),
	.B0 (n_923),
	.A1 (n_868),
	.A0 (n_857) );
   AOI21X1 i_609 ( .Y (n_1011),
	.B0 (n_924),
	.A1 (n_878),
	.A0 (n_869) );
   AOI21X1 i_611 ( .Y (n_1013),
	.B0 (n_925),
	.A1 (n_879),
	.A0 (n_886) );
   AOI21X1 i_613 ( .Y (n_1015),
	.B0 (n_926),
	.A1 (n_892),
	.A0 (n_887) );
   AOI21X1 i_615 ( .Y (n_1017),
	.B0 (n_927),
	.A1 (n_893),
	.A0 (n_896) );
   AOI21X1 i_617 ( .Y (n_1019),
	.B0 (n_928),
	.A1 (n_897),
	.A0 (n_898) );
   AOI31X1 i_619 ( .Y (n_1021),
	.B0 (n_929),
	.A2 (n_899),
	.A1 (a[15]),
	.A0 (b[15]) );
   NOR2X1 i_654 ( .Y (n_1056),
	.B (n_901),
	.A (n_902) );
   NOR2X1 i_655 ( .Y (n_1057),
	.B (n_902),
	.A (n_903) );
   NOR2X1 i_656 ( .Y (n_1058),
	.B (n_903),
	.A (n_904) );
   XNOR2X1 i_893 ( .Y (y[2]),
	.B (n_931),
	.A (n_965) );
   NOR2X1 i_657 ( .Y (n_1059),
	.B (n_904),
	.A (n_905) );
   NOR2X1 i_658 ( .Y (n_1060),
	.B (n_905),
	.A (n_906) );
   NOR2X1 i_659 ( .Y (n_1061),
	.B (n_906),
	.A (n_907) );
   AOI21X1 i_894 ( .Y (y[3]),
	.B0 (n_5393),
	.A1 (n_1025),
	.A0 (n_967) );
   NOR2X1 i_6310 ( .Y (n_5393),
	.B (n_1025),
	.A (n_967) );
   NOR2X1 i_660 ( .Y (n_1062),
	.B (n_907),
	.A (n_908) );
   NOR2X1 i_661 ( .Y (n_1063),
	.B (n_908),
	.A (n_909) );
   NOR2X1 i_662 ( .Y (n_1064),
	.B (n_909),
	.A (n_910) );
   XNOR2X1 i_895 ( .Y (y[4]),
	.B (n_1086),
	.A (n_969) );
   NOR2X1 i_663 ( .Y (n_1065),
	.B (n_910),
	.A (n_911) );
   NOR2X1 i_664 ( .Y (n_1066),
	.B (n_911),
	.A (n_912) );
   NOR2X1 i_665 ( .Y (n_1067),
	.B (n_912),
	.A (n_913) );
   XNOR2X1 i_896 ( .Y (y[5]),
	.B (n_1087),
	.A (n_971) );
   NOR2X1 i_666 ( .Y (n_1068),
	.B (n_913),
	.A (n_914) );
   NOR2X1 i_667 ( .Y (n_1069),
	.B (n_914),
	.A (n_915) );
   NOR2X1 i_668 ( .Y (n_1070),
	.B (n_915),
	.A (n_916) );
   AOI21X1 i_897 ( .Y (y[6]),
	.B0 (n_5408),
	.A1 (n_1148),
	.A0 (n_973) );
   NOR2X1 i_6325 ( .Y (n_5408),
	.B (n_1148),
	.A (n_973) );
   NOR2X1 i_669 ( .Y (n_1071),
	.B (n_916),
	.A (n_917) );
   NOR2X1 i_670 ( .Y (n_1072),
	.B (n_917),
	.A (n_918) );
   NOR2X1 i_671 ( .Y (n_1073),
	.B (n_918),
	.A (n_919) );
   AOI21X1 i_898 ( .Y (y[7]),
	.B0 (n_5413),
	.A1 (n_1149),
	.A0 (n_975) );
   NOR2X1 i_6330 ( .Y (n_5413),
	.B (n_1149),
	.A (n_975) );
   NOR2X1 i_672 ( .Y (n_1074),
	.B (n_919),
	.A (n_920) );
   NOR2X1 i_673 ( .Y (n_1075),
	.B (n_920),
	.A (n_921) );
   NOR2X1 i_674 ( .Y (n_1076),
	.B (n_921),
	.A (n_922) );
   AOI21X1 i_899 ( .Y (y[8]),
	.B0 (n_5418),
	.A1 (n_1150),
	.A0 (n_977) );
   NOR2X1 i_6335 ( .Y (n_5418),
	.B (n_1150),
	.A (n_977) );
   NOR2X1 i_675 ( .Y (n_1077),
	.B (n_922),
	.A (n_923) );
   NOR2X1 i_676 ( .Y (n_1078),
	.B (n_923),
	.A (n_924) );
   NOR2X1 i_677 ( .Y (n_1079),
	.B (n_924),
	.A (n_925) );
   AOI21X1 i_900 ( .Y (y[9]),
	.B0 (n_5423),
	.A1 (n_1151),
	.A0 (n_979) );
   NOR2X1 i_6340 ( .Y (n_5423),
	.B (n_1151),
	.A (n_979) );
   NOR2X1 i_678 ( .Y (n_1080),
	.B (n_925),
	.A (n_926) );
   NOR2X1 i_679 ( .Y (n_1081),
	.B (n_926),
	.A (n_927) );
   NOR2X1 i_680 ( .Y (n_1082),
	.B (n_927),
	.A (n_928) );
   XNOR2X1 i_901 ( .Y (y[10]),
	.B (n_1212),
	.A (n_981) );
   NOR2X1 i_681 ( .Y (n_1083),
	.B (n_928),
	.A (n_929) );
   NAND2X1 i_716 ( .Y (n_1118),
	.B (n_1056),
	.A (n_1058) );
   NAND2X1 i_717 ( .Y (n_1119),
	.B (n_1057),
	.A (n_1059) );
   XNOR2X1 i_902 ( .Y (y[11]),
	.B (n_1213),
	.A (n_983) );
   NAND2X1 i_718 ( .Y (n_1120),
	.B (n_1058),
	.A (n_1060) );
   NAND2X1 i_719 ( .Y (n_1121),
	.B (n_1059),
	.A (n_1061) );
   NAND2X1 i_720 ( .Y (n_1122),
	.B (n_1060),
	.A (n_1062) );
   XNOR2X1 i_903 ( .Y (y[12]),
	.B (n_1214),
	.A (n_985) );
   NAND2X1 i_721 ( .Y (n_1123),
	.B (n_1061),
	.A (n_1063) );
   NAND2X1 i_722 ( .Y (n_1124),
	.B (n_1062),
	.A (n_1064) );
   NAND2X1 i_723 ( .Y (n_1125),
	.B (n_1063),
	.A (n_1065) );
   XNOR2X1 i_904 ( .Y (y[13]),
	.B (n_1215),
	.A (n_987) );
   NAND2X1 i_724 ( .Y (n_1126),
	.B (n_1064),
	.A (n_1066) );
   NAND2X1 i_725 ( .Y (n_1127),
	.B (n_1065),
	.A (n_1067) );
   NAND2X1 i_726 ( .Y (n_1128),
	.B (n_1066),
	.A (n_1068) );
   XNOR2X1 i_905 ( .Y (y[14]),
	.B (n_1216),
	.A (n_989) );
   NAND2X1 i_727 ( .Y (n_1129),
	.B (n_1067),
	.A (n_1069) );
   NAND2X1 i_728 ( .Y (n_1130),
	.B (n_1068),
	.A (n_1070) );
   NAND2X1 i_729 ( .Y (n_1131),
	.B (n_1069),
	.A (n_1071) );
   XNOR2X1 i_906 ( .Y (y[15]),
	.B (n_1217),
	.A (n_991) );
   NAND2X1 i_730 ( .Y (n_1132),
	.B (n_1070),
	.A (n_1072) );
   NAND2X1 i_731 ( .Y (n_1133),
	.B (n_1071),
	.A (n_1073) );
   NAND2X1 i_732 ( .Y (n_1134),
	.B (n_1072),
	.A (n_1074) );
   XNOR2X1 i_907 ( .Y (y[16]),
	.B (n_1218),
	.A (n_993) );
   NAND2X1 i_733 ( .Y (n_1135),
	.B (n_1073),
	.A (n_1075) );
   NAND2X1 i_734 ( .Y (n_1136),
	.B (n_1074),
	.A (n_1076) );
   NAND2X1 i_735 ( .Y (n_1137),
	.B (n_1075),
	.A (n_1077) );
   XNOR2X1 i_908 ( .Y (y[17]),
	.B (n_1219),
	.A (n_995) );
   NAND2X1 i_736 ( .Y (n_1138),
	.B (n_1076),
	.A (n_1078) );
   NAND2X1 i_737 ( .Y (n_1139),
	.B (n_1077),
	.A (n_1079) );
   NAND2X1 i_738 ( .Y (n_1140),
	.B (n_1078),
	.A (n_1080) );
   AOI21X1 i_909 ( .Y (y[18]),
	.B0 (n_5468),
	.A1 (n_1280),
	.A0 (n_997) );
   NOR2X1 i_6385 ( .Y (n_5468),
	.B (n_1280),
	.A (n_997) );
   NAND2X1 i_739 ( .Y (n_1141),
	.B (n_1079),
	.A (n_1081) );
   NAND2X1 i_740 ( .Y (n_1142),
	.B (n_1080),
	.A (n_1082) );
   NAND2X1 i_741 ( .Y (n_1143),
	.B (n_1081),
	.A (n_1083) );
   AOI21X1 i_910 ( .Y (y[19]),
	.B0 (n_5473),
	.A1 (n_1281),
	.A0 (n_999) );
   NOR2X1 i_6390 ( .Y (n_5473),
	.B (n_1281),
	.A (n_999) );
   NOR2X1 i_780 ( .Y (n_1182),
	.B (n_1118),
	.A (n_1122) );
   NOR2X1 i_781 ( .Y (n_1183),
	.B (n_1119),
	.A (n_1123) );
   NOR2X1 i_782 ( .Y (n_1184),
	.B (n_1120),
	.A (n_1124) );
   AOI21X1 i_911 ( .Y (y[20]),
	.B0 (n_5478),
	.A1 (n_1282),
	.A0 (n_1001) );
   NOR2X1 i_6395 ( .Y (n_5478),
	.B (n_1282),
	.A (n_1001) );
   NOR2X1 i_783 ( .Y (n_1185),
	.B (n_1121),
	.A (n_1125) );
   NOR2X1 i_784 ( .Y (n_1186),
	.B (n_1122),
	.A (n_1126) );
   NOR2X1 i_785 ( .Y (n_1187),
	.B (n_1123),
	.A (n_1127) );
   AOI21X1 i_912 ( .Y (y[21]),
	.B0 (n_5483),
	.A1 (n_1283),
	.A0 (n_1003) );
   NOR2X1 i_6400 ( .Y (n_5483),
	.B (n_1283),
	.A (n_1003) );
   NOR2X1 i_786 ( .Y (n_1188),
	.B (n_1124),
	.A (n_1128) );
   NOR2X1 i_787 ( .Y (n_1189),
	.B (n_1125),
	.A (n_1129) );
   NOR2X1 i_788 ( .Y (n_1190),
	.B (n_1126),
	.A (n_1130) );
   AOI21X1 i_913 ( .Y (y[22]),
	.B0 (n_5488),
	.A1 (n_1284),
	.A0 (n_1005) );
   NOR2X1 i_6405 ( .Y (n_5488),
	.B (n_1284),
	.A (n_1005) );
   NOR2X1 i_789 ( .Y (n_1191),
	.B (n_1127),
	.A (n_1131) );
   NOR2X1 i_790 ( .Y (n_1192),
	.B (n_1128),
	.A (n_1132) );
   NOR2X1 i_791 ( .Y (n_1193),
	.B (n_1129),
	.A (n_1133) );
   AOI21X1 i_914 ( .Y (y[23]),
	.B0 (n_5493),
	.A1 (n_1285),
	.A0 (n_1007) );
   NOR2X1 i_6410 ( .Y (n_5493),
	.B (n_1285),
	.A (n_1007) );
   NOR2X1 i_792 ( .Y (n_1194),
	.B (n_1130),
	.A (n_1134) );
   NOR2X1 i_793 ( .Y (n_1195),
	.B (n_1131),
	.A (n_1135) );
   NOR2X1 i_794 ( .Y (n_1196),
	.B (n_1132),
	.A (n_1136) );
   AOI21X1 i_915 ( .Y (y[24]),
	.B0 (n_5498),
	.A1 (n_1286),
	.A0 (n_1009) );
   NOR2X1 i_6415 ( .Y (n_5498),
	.B (n_1286),
	.A (n_1009) );
   NOR2X1 i_795 ( .Y (n_1197),
	.B (n_1133),
	.A (n_1137) );
   NOR2X1 i_796 ( .Y (n_1198),
	.B (n_1134),
	.A (n_1138) );
   NOR2X1 i_797 ( .Y (n_1199),
	.B (n_1135),
	.A (n_1139) );
   AOI21X1 i_916 ( .Y (y[25]),
	.B0 (n_5503),
	.A1 (n_1287),
	.A0 (n_1011) );
   NOR2X1 i_6420 ( .Y (n_5503),
	.B (n_1287),
	.A (n_1011) );
   NOR2X1 i_798 ( .Y (n_1200),
	.B (n_1136),
	.A (n_1140) );
   NOR2X1 i_799 ( .Y (n_1201),
	.B (n_1137),
	.A (n_1141) );
   NOR2X1 i_800 ( .Y (n_1202),
	.B (n_1138),
	.A (n_1142) );
   AOI21X1 i_917 ( .Y (y[26]),
	.B0 (n_5508),
	.A1 (n_1288),
	.A0 (n_1013) );
   NOR2X1 i_6425 ( .Y (n_5508),
	.B (n_1288),
	.A (n_1013) );
   NOR2X1 i_801 ( .Y (n_1203),
	.B (n_1139),
	.A (n_1143) );
   NAND2X1 i_848 ( .Y (n_1250),
	.B (n_1190),
	.A (n_1182) );
   NAND2X1 i_849 ( .Y (n_1251),
	.B (n_1191),
	.A (n_1183) );
   AOI21X1 i_918 ( .Y (y[27]),
	.B0 (n_5513),
	.A1 (n_1289),
	.A0 (n_1015) );
   NOR2X1 i_6430 ( .Y (n_5513),
	.B (n_1289),
	.A (n_1015) );
   NAND2X1 i_850 ( .Y (n_1252),
	.B (n_1192),
	.A (n_1184) );
   NAND2X1 i_851 ( .Y (n_1253),
	.B (n_1193),
	.A (n_1185) );
   NAND2X1 i_852 ( .Y (n_1254),
	.B (n_1194),
	.A (n_1186) );
   AOI21X1 i_919 ( .Y (y[28]),
	.B0 (n_5518),
	.A1 (n_1290),
	.A0 (n_1017) );
   NOR2X1 i_6435 ( .Y (n_5518),
	.B (n_1290),
	.A (n_1017) );
   NAND2X1 i_853 ( .Y (n_1255),
	.B (n_1187),
	.A (n_1195) );
   NAND2X1 i_854 ( .Y (n_1256),
	.B (n_1196),
	.A (n_1188) );
   NAND2X1 i_855 ( .Y (n_1257),
	.B (n_1197),
	.A (n_1189) );
   AOI21X1 i_920 ( .Y (y[29]),
	.B0 (n_5523),
	.A1 (n_1291),
	.A0 (n_1019) );
   NOR2X1 i_6440 ( .Y (n_5523),
	.B (n_1291),
	.A (n_1019) );
   NAND2X1 i_856 ( .Y (n_1258),
	.B (n_1198),
	.A (n_1190) );
   NAND2X1 i_857 ( .Y (n_1259),
	.B (n_1199),
	.A (n_1191) );
   NAND4BXL i_858 ( .Y (n_1260),
	.D (n_1192),
	.C (n_1078),
	.B (n_1080),
	.AN (n_1136) );
   AOI21X1 i_921 ( .Y (y[30]),
	.B0 (n_5528),
	.A1 (n_1292),
	.A0 (n_1021) );
   NOR2X1 i_6445 ( .Y (n_5528),
	.B (n_1292),
	.A (n_1021) );
   NAND4BXL i_859 ( .Y (n_1261),
	.D (n_1193),
	.C (n_1079),
	.B (n_1081),
	.AN (n_1137) );
   NAND4BXL i_860 ( .Y (n_1262),
	.D (n_1194),
	.C (n_1080),
	.B (n_1082),
	.AN (n_1138) );
   NAND2X1 i_861 ( .Y (n_1263),
	.B (n_1195),
	.A (n_1203) );
   INVX1 i_6930 ( .Y (n_1211),
	.A (n_1151) );
   INVX1 i_6931 ( .Y (n_1210),
	.A (n_1150) );
   INVX1 i_6932 ( .Y (n_1209),
	.A (n_1149) );
   INVX1 i_6933 ( .Y (n_1208),
	.A (n_1148) );
   INVX1 i_6934 ( .Y (n_1085),
	.A (n_1025) );
   INVX1 i_6935 ( .Y (n_1147),
	.A (n_1087) );
   INVX1 i_6936 ( .Y (n_1146),
	.A (n_1086) );
   INVX1 i_6937 ( .Y (n_931),
	.A (n_1024) );
   ADDHX1 i_288 ( .S (n_480),
	.CO (n_481),
	.B (n_448),
	.A (n_466) );
   ADDHX1 i_289 ( .S (n_482),
	.CO (n_483),
	.B (n_449),
	.A (n_467) );
   ADDFHX1 i_290 ( .S (n_484),
	.CO (n_485),
	.CI (n_481),
	.B (n_413),
	.A (n_431) );
   ADDHX1 i_291 ( .S (n_486),
	.CO (n_487),
	.B (n_450),
	.A (n_468) );
   ADDFHX1 i_292 ( .S (n_488),
	.CO (n_489),
	.CI (n_396),
	.B (n_414),
	.A (n_432) );
   ADDFHX1 i_293 ( .S (n_490),
	.CO (n_491),
	.CI (n_488),
	.B (n_486),
	.A (n_483) );
   ADDHX1 i_294 ( .S (n_492),
	.CO (n_493),
	.B (n_451),
	.A (n_469) );
   ADDFHX1 i_295 ( .S (n_494),
	.CO (n_495),
	.CI (n_397),
	.B (n_415),
	.A (n_433) );
   ADDFHX1 i_296 ( .S (n_496),
	.CO (n_497),
	.CI (n_489),
	.B (n_487),
	.A (n_379) );
   ADDFHX1 i_297 ( .S (n_498),
	.CO (n_499),
	.CI (n_491),
	.B (n_494),
	.A (n_492) );
   ADDHX1 i_298 ( .S (n_500),
	.CO (n_501),
	.B (n_452),
	.A (n_470) );
   ADDFHX1 i_299 ( .S (n_502),
	.CO (n_503),
	.CI (n_398),
	.B (n_416),
	.A (n_434) );
   ADDFHX1 i_300 ( .S (n_504),
	.CO (n_505),
	.CI (n_493),
	.B (n_362),
	.A (n_380) );
   ADDFHX1 i_301 ( .S (n_506),
	.CO (n_507),
	.CI (n_502),
	.B (n_500),
	.A (n_495) );
   ADDFHX1 i_302 ( .S (n_508),
	.CO (n_509),
	.CI (n_506),
	.B (n_504),
	.A (n_497) );
   ADDHX1 i_303 ( .S (n_510),
	.CO (n_511),
	.B (n_453),
	.A (n_471) );
   ADDFHX1 i_304 ( .S (n_512),
	.CO (n_513),
	.CI (n_399),
	.B (n_417),
	.A (n_435) );
   ADDFHX1 i_305 ( .S (n_514),
	.CO (n_515),
	.CI (n_345),
	.B (n_363),
	.A (n_381) );
   ADDFHX1 i_306 ( .S (n_516),
	.CO (n_517),
	.CI (n_510),
	.B (n_503),
	.A (n_501) );
   ADDFHX1 i_307 ( .S (n_518),
	.CO (n_519),
	.CI (n_505),
	.B (n_514),
	.A (n_512) );
   ADDFHX1 i_308 ( .S (n_520),
	.CO (n_521),
	.CI (n_509),
	.B (n_516),
	.A (n_507) );
   ADDHX1 i_309 ( .S (n_522),
	.CO (n_523),
	.B (n_454),
	.A (n_472) );
   ADDFHX1 i_310 ( .S (n_524),
	.CO (n_525),
	.CI (n_400),
	.B (n_418),
	.A (n_436) );
   ADDFHX1 i_311 ( .S (n_526),
	.CO (n_527),
	.CI (n_346),
	.B (n_364),
	.A (n_382) );
   ADDFHX1 i_312 ( .S (n_528),
	.CO (n_529),
	.CI (n_513),
	.B (n_511),
	.A (n_328) );
   ADDFHX1 i_313 ( .S (n_530),
	.CO (n_531),
	.CI (n_524),
	.B (n_522),
	.A (n_515) );
   ADDFHX1 i_314 ( .S (n_532),
	.CO (n_533),
	.CI (n_528),
	.B (n_517),
	.A (n_526) );
   ADDFHX1 i_315 ( .S (n_534),
	.CO (n_535),
	.CI (n_532),
	.B (n_519),
	.A (n_530) );
   ADDHX1 i_316 ( .S (n_536),
	.CO (n_537),
	.B (n_455),
	.A (n_473) );
   ADDFHX1 i_317 ( .S (n_538),
	.CO (n_539),
	.CI (n_401),
	.B (n_419),
	.A (n_437) );
   ADDFHX1 i_318 ( .S (n_540),
	.CO (n_541),
	.CI (n_347),
	.B (n_365),
	.A (n_383) );
   ADDFHX1 i_319 ( .S (n_542),
	.CO (n_543),
	.CI (n_523),
	.B (n_311),
	.A (n_329) );
   ADDFHX1 i_320 ( .S (n_544),
	.CO (n_545),
	.CI (n_536),
	.B (n_527),
	.A (n_525) );
   ADDFHX1 i_321 ( .S (n_546),
	.CO (n_547),
	.CI (n_529),
	.B (n_540),
	.A (n_538) );
   ADDFHX1 i_322 ( .S (n_548),
	.CO (n_549),
	.CI (n_544),
	.B (n_542),
	.A (n_531) );
   ADDFHX1 i_323 ( .S (n_550),
	.CO (n_551),
	.CI (n_548),
	.B (n_546),
	.A (n_533) );
   ADDHX1 i_324 ( .S (n_552),
	.CO (n_553),
	.B (n_456),
	.A (n_474) );
   ADDFHX1 i_325 ( .S (n_554),
	.CO (n_555),
	.CI (n_402),
	.B (n_420),
	.A (n_438) );
   ADDFHX1 i_326 ( .S (n_556),
	.CO (n_557),
	.CI (n_348),
	.B (n_366),
	.A (n_384) );
   ADDFHX1 i_327 ( .S (n_558),
	.CO (n_559),
	.CI (n_294),
	.B (n_312),
	.A (n_330) );
   ADDFHX1 i_328 ( .S (n_560),
	.CO (n_561),
	.CI (n_541),
	.B (n_539),
	.A (n_537) );
   ADDFHX1 i_329 ( .S (n_562),
	.CO (n_563),
	.CI (n_556),
	.B (n_554),
	.A (n_552) );
   ADDFHX1 i_330 ( .S (n_564),
	.CO (n_565),
	.CI (n_545),
	.B (n_543),
	.A (n_558) );
   ADDFHX1 i_331 ( .S (n_566),
	.CO (n_567),
	.CI (n_547),
	.B (n_562),
	.A (n_560) );
   ADDFHX1 i_332 ( .S (n_568),
	.CO (n_569),
	.CI (n_551),
	.B (n_564),
	.A (n_549) );
   ADDHX1 i_333 ( .S (n_570),
	.CO (n_571),
	.B (n_457),
	.A (n_475) );
   ADDFHX1 i_334 ( .S (n_572),
	.CO (n_573),
	.CI (n_403),
	.B (n_421),
	.A (n_439) );
   ADDFHX1 i_335 ( .S (n_574),
	.CO (n_575),
	.CI (n_349),
	.B (n_367),
	.A (n_385) );
   ADDFHX1 i_336 ( .S (n_576),
	.CO (n_577),
	.CI (n_295),
	.B (n_313),
	.A (n_331) );
   ADDFHX1 i_337 ( .S (n_578),
	.CO (n_579),
	.CI (n_555),
	.B (n_553),
	.A (n_277) );
   ADDFHX1 i_338 ( .S (n_580),
	.CO (n_581),
	.CI (n_570),
	.B (n_559),
	.A (n_557) );
   ADDFHX1 i_339 ( .S (n_582),
	.CO (n_583),
	.CI (n_576),
	.B (n_574),
	.A (n_572) );
   ADDFHX1 i_340 ( .S (n_584),
	.CO (n_585),
	.CI (n_578),
	.B (n_563),
	.A (n_561) );
   ADDFHX1 i_341 ( .S (n_586),
	.CO (n_587),
	.CI (n_565),
	.B (n_582),
	.A (n_580) );
   ADDFHX1 i_342 ( .S (n_588),
	.CO (n_589),
	.CI (n_586),
	.B (n_567),
	.A (n_584) );
   ADDHX1 i_343 ( .S (n_590),
	.CO (n_591),
	.B (n_458),
	.A (n_476) );
   ADDFHX1 i_344 ( .S (n_592),
	.CO (n_593),
	.CI (n_404),
	.B (n_422),
	.A (n_440) );
   ADDFHX1 i_345 ( .S (n_594),
	.CO (n_595),
	.CI (n_350),
	.B (n_368),
	.A (n_386) );
   ADDFHX1 i_346 ( .S (n_596),
	.CO (n_597),
	.CI (n_296),
	.B (n_314),
	.A (n_332) );
   ADDFHX1 i_347 ( .S (n_598),
	.CO (n_599),
	.CI (n_571),
	.B (n_260),
	.A (n_278) );
   ADDFHX1 i_348 ( .S (n_600),
	.CO (n_601),
	.CI (n_577),
	.B (n_575),
	.A (n_573) );
   ADDFHX1 i_349 ( .S (n_602),
	.CO (n_603),
	.CI (n_594),
	.B (n_592),
	.A (n_590) );
   ADDFHX1 i_350 ( .S (n_604),
	.CO (n_605),
	.CI (n_581),
	.B (n_579),
	.A (n_596) );
   ADDFHX1 i_351 ( .S (n_606),
	.CO (n_607),
	.CI (n_600),
	.B (n_598),
	.A (n_583) );
   ADDFHX1 i_352 ( .S (n_608),
	.CO (n_609),
	.CI (n_604),
	.B (n_585),
	.A (n_602) );
   ADDFHX1 i_353 ( .S (n_610),
	.CO (n_611),
	.CI (n_608),
	.B (n_587),
	.A (n_606) );
   ADDHX1 i_354 ( .S (n_612),
	.CO (n_613),
	.B (n_459),
	.A (n_477) );
   ADDFHX1 i_355 ( .S (n_614),
	.CO (n_615),
	.CI (n_405),
	.B (n_423),
	.A (n_441) );
   ADDFHX1 i_356 ( .S (n_616),
	.CO (n_617),
	.CI (n_351),
	.B (n_369),
	.A (n_387) );
   ADDFHX1 i_357 ( .S (n_618),
	.CO (n_619),
	.CI (n_297),
	.B (n_315),
	.A (n_333) );
   ADDFHX1 i_358 ( .S (n_620),
	.CO (n_621),
	.CI (n_243),
	.B (n_261),
	.A (n_279) );
   ADDFHX1 i_359 ( .S (n_622),
	.CO (n_623),
	.CI (n_595),
	.B (n_593),
	.A (n_591) );
   ADDFHX1 i_360 ( .S (n_624),
	.CO (n_625),
	.CI (n_614),
	.B (n_612),
	.A (n_597) );
   ADDFHX1 i_361 ( .S (n_626),
	.CO (n_627),
	.CI (n_620),
	.B (n_618),
	.A (n_616) );
   ADDFHX1 i_362 ( .S (n_628),
	.CO (n_629),
	.CI (n_603),
	.B (n_601),
	.A (n_599) );
   ADDFHX1 i_363 ( .S (n_630),
	.CO (n_631),
	.CI (n_626),
	.B (n_624),
	.A (n_622) );
   ADDFHX1 i_364 ( .S (n_632),
	.CO (n_633),
	.CI (n_628),
	.B (n_607),
	.A (n_605) );
   ADDFHX1 i_365 ( .S (n_634),
	.CO (n_635),
	.CI (n_632),
	.B (n_609),
	.A (n_630) );
   ADDHX1 i_366 ( .S (n_636),
	.CO (n_637),
	.B (n_460),
	.A (n_478) );
   ADDFHX1 i_367 ( .S (n_638),
	.CO (n_639),
	.CI (n_406),
	.B (n_424),
	.A (n_442) );
   ADDFHX1 i_368 ( .S (n_640),
	.CO (n_641),
	.CI (n_352),
	.B (n_370),
	.A (n_388) );
   ADDFHX1 i_369 ( .S (n_642),
	.CO (n_643),
	.CI (n_298),
	.B (n_316),
	.A (n_334) );
   ADDFHX1 i_370 ( .S (n_644),
	.CO (n_645),
	.CI (n_244),
	.B (n_262),
	.A (n_280) );
   ADDFHX1 i_371 ( .S (n_646),
	.CO (n_647),
	.CI (n_615),
	.B (n_613),
	.A (n_226) );
   ADDFHX1 i_372 ( .S (n_648),
	.CO (n_649),
	.CI (n_621),
	.B (n_619),
	.A (n_617) );
   ADDFHX1 i_373 ( .S (n_650),
	.CO (n_651),
	.CI (n_640),
	.B (n_638),
	.A (n_636) );
   ADDFHX1 i_374 ( .S (n_652),
	.CO (n_653),
	.CI (n_623),
	.B (n_644),
	.A (n_642) );
   ADDFHX1 i_375 ( .S (n_654),
	.CO (n_655),
	.CI (n_646),
	.B (n_627),
	.A (n_625) );
   ADDFHX1 i_376 ( .S (n_656),
	.CO (n_657),
	.CI (n_629),
	.B (n_650),
	.A (n_648) );
   ADDFHX1 i_377 ( .S (n_658),
	.CO (n_659),
	.CI (n_654),
	.B (n_652),
	.A (n_631) );
   ADDFHX1 i_378 ( .S (n_660),
	.CO (n_661),
	.CI (n_658),
	.B (n_656),
	.A (n_633) );
   ADDHX1 i_379 ( .S (n_662),
	.CO (n_663),
	.B (n_461),
	.A (n_479) );
   ADDFHX1 i_380 ( .S (n_664),
	.CO (n_665),
	.CI (n_407),
	.B (n_425),
	.A (n_443) );
   ADDFHX1 i_381 ( .S (n_666),
	.CO (n_667),
	.CI (n_353),
	.B (n_371),
	.A (n_389) );
   ADDFHX1 i_382 ( .S (n_668),
	.CO (n_669),
	.CI (n_299),
	.B (n_317),
	.A (n_335) );
   ADDFHX1 i_383 ( .S (n_670),
	.CO (n_671),
	.CI (n_245),
	.B (n_263),
	.A (n_281) );
   ADDFHX1 i_384 ( .S (n_672),
	.CO (n_673),
	.CI (n_637),
	.B (n_209),
	.A (n_227) );
   ADDFHX1 i_385 ( .S (n_674),
	.CO (n_675),
	.CI (n_643),
	.B (n_641),
	.A (n_639) );
   ADDFHX1 i_386 ( .S (n_676),
	.CO (n_677),
	.CI (n_664),
	.B (n_662),
	.A (n_645) );
   ADDFHX1 i_387 ( .S (n_678),
	.CO (n_679),
	.CI (n_670),
	.B (n_668),
	.A (n_666) );
   ADDFHX1 i_388 ( .S (n_680),
	.CO (n_681),
	.CI (n_651),
	.B (n_649),
	.A (n_647) );
   ADDFHX1 i_389 ( .S (n_682),
	.CO (n_683),
	.CI (n_676),
	.B (n_674),
	.A (n_672) );
   ADDFHX1 i_390 ( .S (n_684),
	.CO (n_685),
	.CI (n_655),
	.B (n_653),
	.A (n_678) );
   ADDFHX1 i_391 ( .S (n_686),
	.CO (n_687),
	.CI (n_657),
	.B (n_682),
	.A (n_680) );
   ADDFHX1 i_392 ( .S (n_688),
	.CO (n_689),
	.CI (n_661),
	.B (n_684),
	.A (n_659) );
   ADDHX1 i_393 ( .S (n_690),
	.CO (n_691),
	.B (n_444),
	.A (n_462) );
   ADDFHX1 i_394 ( .S (n_692),
	.CO (n_693),
	.CI (n_390),
	.B (n_408),
	.A (n_426) );
   ADDFHX1 i_395 ( .S (n_694),
	.CO (n_695),
	.CI (n_336),
	.B (n_354),
	.A (n_372) );
   ADDFHX1 i_396 ( .S (n_696),
	.CO (n_697),
	.CI (n_282),
	.B (n_300),
	.A (n_318) );
   ADDFHX1 i_397 ( .S (n_698),
	.CO (n_699),
	.CI (n_228),
	.B (n_246),
	.A (n_264) );
   ADDFHX1 i_398 ( .S (n_700),
	.CO (n_701),
	.CI (n_665),
	.B (n_663),
	.A (n_210) );
   ADDFHX1 i_399 ( .S (n_702),
	.CO (n_703),
	.CI (n_671),
	.B (n_669),
	.A (n_667) );
   ADDFHX1 i_400 ( .S (n_704),
	.CO (n_705),
	.CI (n_694),
	.B (n_692),
	.A (n_690) );
   ADDFHX1 i_401 ( .S (n_706),
	.CO (n_707),
	.CI (n_673),
	.B (n_698),
	.A (n_696) );
   ADDFHX1 i_402 ( .S (n_708),
	.CO (n_709),
	.CI (n_679),
	.B (n_677),
	.A (n_675) );
   ADDFHX1 i_403 ( .S (n_710),
	.CO (n_711),
	.CI (n_704),
	.B (n_702),
	.A (n_700) );
   ADDFHX1 i_404 ( .S (n_712),
	.CO (n_713),
	.CI (n_706),
	.B (n_683),
	.A (n_681) );
   ADDFHX1 i_405 ( .S (n_714),
	.CO (n_715),
	.CI (n_685),
	.B (n_710),
	.A (n_708) );
   ADDFHX1 i_406 ( .S (n_716),
	.CO (n_717),
	.CI (n_714),
	.B (n_687),
	.A (n_712) );
   ADDFHX1 i_407 ( .S (n_718),
	.CO (n_719),
	.CI (n_409),
	.B (n_427),
	.A (n_445) );
   ADDFHX1 i_408 ( .S (n_720),
	.CO (n_721),
	.CI (n_355),
	.B (n_373),
	.A (n_391) );
   ADDFHX1 i_409 ( .S (n_722),
	.CO (n_723),
	.CI (n_301),
	.B (n_319),
	.A (n_337) );
   ADDFHX1 i_410 ( .S (n_724),
	.CO (n_725),
	.CI (n_247),
	.B (n_265),
	.A (n_283) );
   ADDFHX1 i_411 ( .S (n_726),
	.CO (n_727),
	.CI (n_691),
	.B (n_211),
	.A (n_229) );
   ADDFHX1 i_412 ( .S (n_728),
	.CO (n_729),
	.CI (n_697),
	.B (n_695),
	.A (n_693) );
   ADDFHX1 i_413 ( .S (n_730),
	.CO (n_731),
	.CI (n_720),
	.B (n_718),
	.A (n_699) );
   ADDFHX1 i_414 ( .S (n_732),
	.CO (n_733),
	.CI (n_701),
	.B (n_724),
	.A (n_722) );
   ADDFHX1 i_415 ( .S (n_734),
	.CO (n_735),
	.CI (n_726),
	.B (n_705),
	.A (n_703) );
   ADDFHX1 i_416 ( .S (n_736),
	.CO (n_737),
	.CI (n_707),
	.B (n_730),
	.A (n_728) );
   ADDFHX1 i_417 ( .S (n_738),
	.CO (n_739),
	.CI (n_732),
	.B (n_711),
	.A (n_709) );
   ADDFHX1 i_418 ( .S (n_740),
	.CO (n_741),
	.CI (n_736),
	.B (n_713),
	.A (n_734) );
   ADDFHX1 i_419 ( .S (n_742),
	.CO (n_743),
	.CI (n_740),
	.B (n_715),
	.A (n_738) );
   ADDFHX1 i_420 ( .S (n_744),
	.CO (n_745),
	.CI (n_392),
	.B (n_410),
	.A (n_428) );
   ADDFHX1 i_421 ( .S (n_746),
	.CO (n_747),
	.CI (n_338),
	.B (n_356),
	.A (n_374) );
   ADDFHX1 i_422 ( .S (n_748),
	.CO (n_749),
	.CI (n_284),
	.B (n_302),
	.A (n_320) );
   ADDFHX1 i_423 ( .S (n_750),
	.CO (n_751),
	.CI (n_230),
	.B (n_248),
	.A (n_266) );
   ADDFHX1 i_424 ( .S (n_752),
	.CO (n_753),
	.CI (n_721),
	.B (n_719),
	.A (n_212) );
   ADDFHX1 i_425 ( .S (n_754),
	.CO (n_755),
	.CI (n_744),
	.B (n_725),
	.A (n_723) );
   ADDFHX1 i_426 ( .S (n_756),
	.CO (n_757),
	.CI (n_750),
	.B (n_748),
	.A (n_746) );
   ADDFHX1 i_427 ( .S (n_758),
	.CO (n_759),
	.CI (n_731),
	.B (n_729),
	.A (n_727) );
   ADDFHX1 i_428 ( .S (n_760),
	.CO (n_761),
	.CI (n_756),
	.B (n_754),
	.A (n_752) );
   ADDFHX1 i_429 ( .S (n_762),
	.CO (n_763),
	.CI (n_758),
	.B (n_735),
	.A (n_733) );
   ADDFHX1 i_430 ( .S (n_764),
	.CO (n_765),
	.CI (n_739),
	.B (n_737),
	.A (n_760) );
   ADDFHX1 i_431 ( .S (n_766),
	.CO (n_767),
	.CI (n_764),
	.B (n_741),
	.A (n_762) );
   ADDFHX1 i_432 ( .S (n_768),
	.CO (n_769),
	.CI (n_375),
	.B (n_393),
	.A (n_411) );
   ADDFHX1 i_433 ( .S (n_770),
	.CO (n_771),
	.CI (n_321),
	.B (n_339),
	.A (n_357) );
   ADDFHX1 i_434 ( .S (n_772),
	.CO (n_773),
	.CI (n_267),
	.B (n_285),
	.A (n_303) );
   ADDFHX1 i_435 ( .S (n_774),
	.CO (n_775),
	.CI (n_213),
	.B (n_231),
	.A (n_249) );
   ADDFHX1 i_436 ( .S (n_776),
	.CO (n_777),
	.CI (n_749),
	.B (n_747),
	.A (n_745) );
   ADDFHX1 i_437 ( .S (n_778),
	.CO (n_779),
	.CI (n_770),
	.B (n_768),
	.A (n_751) );
   ADDFHX1 i_438 ( .S (n_780),
	.CO (n_781),
	.CI (n_753),
	.B (n_774),
	.A (n_772) );
   ADDFHX1 i_439 ( .S (n_782),
	.CO (n_783),
	.CI (n_776),
	.B (n_757),
	.A (n_755) );
   ADDFHX1 i_440 ( .S (n_784),
	.CO (n_785),
	.CI (n_761),
	.B (n_759),
	.A (n_778) );
   ADDFHX1 i_441 ( .S (n_786),
	.CO (n_787),
	.CI (n_763),
	.B (n_782),
	.A (n_780) );
   ADDFHX1 i_442 ( .S (n_788),
	.CO (n_789),
	.CI (n_786),
	.B (n_765),
	.A (n_784) );
   ADDFHX1 i_443 ( .S (n_790),
	.CO (n_791),
	.CI (n_358),
	.B (n_376),
	.A (n_394) );
   ADDFHX1 i_444 ( .S (n_792),
	.CO (n_793),
	.CI (n_304),
	.B (n_322),
	.A (n_340) );
   ADDFHX1 i_445 ( .S (n_794),
	.CO (n_795),
	.CI (n_250),
	.B (n_268),
	.A (n_286) );
   ADDFHX1 i_446 ( .S (n_796),
	.CO (n_797),
	.CI (n_769),
	.B (n_214),
	.A (n_232) );
   ADDFHX1 i_447 ( .S (n_798),
	.CO (n_799),
	.CI (n_775),
	.B (n_773),
	.A (n_771) );
   ADDFHX1 i_448 ( .S (n_800),
	.CO (n_801),
	.CI (n_794),
	.B (n_792),
	.A (n_790) );
   ADDFHX1 i_449 ( .S (n_802),
	.CO (n_803),
	.CI (n_796),
	.B (n_779),
	.A (n_777) );
   ADDFHX1 i_450 ( .S (n_804),
	.CO (n_805),
	.CI (n_781),
	.B (n_800),
	.A (n_798) );
   ADDFHX1 i_451 ( .S (n_806),
	.CO (n_807),
	.CI (n_785),
	.B (n_802),
	.A (n_783) );
   ADDFHX1 i_452 ( .S (n_808),
	.CO (n_809),
	.CI (n_806),
	.B (n_787),
	.A (n_804) );
   ADDFHX1 i_453 ( .S (n_810),
	.CO (n_811),
	.CI (n_341),
	.B (n_359),
	.A (n_377) );
   ADDFHX1 i_454 ( .S (n_812),
	.CO (n_813),
	.CI (n_287),
	.B (n_305),
	.A (n_323) );
   ADDFHX1 i_455 ( .S (n_814),
	.CO (n_815),
	.CI (n_233),
	.B (n_251),
	.A (n_269) );
   ADDFHX1 i_456 ( .S (n_816),
	.CO (n_817),
	.CI (n_793),
	.B (n_791),
	.A (n_215) );
   ADDFHX1 i_457 ( .S (n_818),
	.CO (n_819),
	.CI (n_812),
	.B (n_810),
	.A (n_795) );
   ADDFHX1 i_458 ( .S (n_820),
	.CO (n_821),
	.CI (n_799),
	.B (n_797),
	.A (n_814) );
   ADDFHX1 i_459 ( .S (n_822),
	.CO (n_823),
	.CI (n_818),
	.B (n_816),
	.A (n_801) );
   ADDFHX1 i_460 ( .S (n_824),
	.CO (n_825),
	.CI (n_822),
	.B (n_820),
	.A (n_803) );
   ADDFHX1 i_461 ( .S (n_826),
	.CO (n_827),
	.CI (n_807),
	.B (n_824),
	.A (n_805) );
   ADDFHX1 i_462 ( .S (n_828),
	.CO (n_829),
	.CI (n_324),
	.B (n_342),
	.A (n_360) );
   ADDFHX1 i_463 ( .S (n_830),
	.CO (n_831),
	.CI (n_270),
	.B (n_288),
	.A (n_306) );
   ADDFHX1 i_464 ( .S (n_832),
	.CO (n_833),
	.CI (n_216),
	.B (n_234),
	.A (n_252) );
   ADDFHX1 i_465 ( .S (n_834),
	.CO (n_835),
	.CI (n_815),
	.B (n_813),
	.A (n_811) );
   ADDFHX1 i_466 ( .S (n_836),
	.CO (n_837),
	.CI (n_832),
	.B (n_830),
	.A (n_828) );
   ADDFHX1 i_467 ( .S (n_838),
	.CO (n_839),
	.CI (n_834),
	.B (n_819),
	.A (n_817) );
   ADDFHX1 i_468 ( .S (n_840),
	.CO (n_841),
	.CI (n_823),
	.B (n_821),
	.A (n_836) );
   ADDFHX1 i_469 ( .S (n_842),
	.CO (n_843),
	.CI (n_840),
	.B (n_825),
	.A (n_838) );
   ADDFHX1 i_470 ( .S (n_844),
	.CO (n_845),
	.CI (n_307),
	.B (n_325),
	.A (n_343) );
   ADDFHX1 i_471 ( .S (n_846),
	.CO (n_847),
	.CI (n_253),
	.B (n_271),
	.A (n_289) );
   ADDFHX1 i_472 ( .S (n_848),
	.CO (n_849),
	.CI (n_829),
	.B (n_217),
	.A (n_235) );
   ADDFHX1 i_473 ( .S (n_850),
	.CO (n_851),
	.CI (n_844),
	.B (n_833),
	.A (n_831) );
   ADDFHX1 i_474 ( .S (n_852),
	.CO (n_853),
	.CI (n_837),
	.B (n_835),
	.A (n_846) );
   ADDFHX1 i_475 ( .S (n_854),
	.CO (n_855),
	.CI (n_839),
	.B (n_850),
	.A (n_848) );
   ADDFHX1 i_476 ( .S (n_856),
	.CO (n_857),
	.CI (n_854),
	.B (n_841),
	.A (n_852) );
   ADDFHX1 i_477 ( .S (n_858),
	.CO (n_859),
	.CI (n_290),
	.B (n_308),
	.A (n_326) );
   ADDFHX1 i_478 ( .S (n_860),
	.CO (n_861),
	.CI (n_236),
	.B (n_254),
	.A (n_272) );
   ADDFHX1 i_479 ( .S (n_862),
	.CO (n_863),
	.CI (n_847),
	.B (n_845),
	.A (n_218) );
   ADDFHX1 i_480 ( .S (n_864),
	.CO (n_865),
	.CI (n_849),
	.B (n_860),
	.A (n_858) );
   ADDFHX1 i_481 ( .S (n_866),
	.CO (n_867),
	.CI (n_853),
	.B (n_862),
	.A (n_851) );
   ADDFHX1 i_482 ( .S (n_868),
	.CO (n_869),
	.CI (n_866),
	.B (n_855),
	.A (n_864) );
   ADDFHX1 i_483 ( .S (n_870),
	.CO (n_871),
	.CI (n_273),
	.B (n_291),
	.A (n_309) );
   ADDFHX1 i_484 ( .S (n_872),
	.CO (n_873),
	.CI (n_219),
	.B (n_237),
	.A (n_255) );
   ADDFHX1 i_485 ( .S (n_874),
	.CO (n_875),
	.CI (n_870),
	.B (n_861),
	.A (n_859) );
   ADDFHX1 i_486 ( .S (n_876),
	.CO (n_877),
	.CI (n_874),
	.B (n_863),
	.A (n_872) );
   ADDFHX1 i_487 ( .S (n_878),
	.CO (n_879),
	.CI (n_867),
	.B (n_876),
	.A (n_865) );
   ADDFHX1 i_488 ( .S (n_880),
	.CO (n_881),
	.CI (n_256),
	.B (n_274),
	.A (n_292) );
   ADDFHX1 i_489 ( .S (n_882),
	.CO (n_883),
	.CI (n_871),
	.B (n_220),
	.A (n_238) );
   ADDFHX1 i_490 ( .S (n_884),
	.CO (n_885),
	.CI (n_875),
	.B (n_880),
	.A (n_873) );
   ADDFHX1 i_491 ( .S (n_886),
	.CO (n_887),
	.CI (n_884),
	.B (n_877),
	.A (n_882) );
   ADDFHX1 i_492 ( .S (n_888),
	.CO (n_889),
	.CI (n_239),
	.B (n_257),
	.A (n_275) );
   ADDFHX1 i_493 ( .S (n_890),
	.CO (n_891),
	.CI (n_888),
	.B (n_881),
	.A (n_221) );
   ADDFHX1 i_494 ( .S (n_892),
	.CO (n_893),
	.CI (n_885),
	.B (n_890),
	.A (n_883) );
   ADDFHX1 i_495 ( .S (n_894),
	.CO (n_895),
	.CI (n_222),
	.B (n_240),
	.A (n_258) );
   ADDFHX1 i_496 ( .S (n_896),
	.CO (n_897),
	.CI (n_891),
	.B (n_894),
	.A (n_889) );
   ADDFHX1 i_497 ( .S (n_898),
	.CO (n_899),
	.CI (n_895),
	.B (n_223),
	.A (n_241) );
   OAI21X1 i_623 ( .Y (n_1025),
	.B0 (n_932),
	.A1 (n_901),
	.A0 (n_931) );
   OAI21X1 i_624 ( .Y (n_1026),
	.B0 (n_933),
	.A1 (n_902),
	.A0 (n_932) );
   OAI21X1 i_625 ( .Y (n_1027),
	.B0 (n_934),
	.A1 (n_903),
	.A0 (n_933) );
   OAI21X1 i_626 ( .Y (n_1028),
	.B0 (n_935),
	.A1 (n_904),
	.A0 (n_934) );
   OAI21X1 i_627 ( .Y (n_1029),
	.B0 (n_936),
	.A1 (n_905),
	.A0 (n_935) );
   OAI21X1 i_628 ( .Y (n_1030),
	.B0 (n_937),
	.A1 (n_906),
	.A0 (n_936) );
   OAI21X1 i_629 ( .Y (n_1031),
	.B0 (n_938),
	.A1 (n_907),
	.A0 (n_937) );
   OAI21X1 i_630 ( .Y (n_1032),
	.B0 (n_939),
	.A1 (n_908),
	.A0 (n_938) );
   OAI21X1 i_631 ( .Y (n_1033),
	.B0 (n_940),
	.A1 (n_909),
	.A0 (n_939) );
   OAI21X1 i_632 ( .Y (n_1034),
	.B0 (n_941),
	.A1 (n_910),
	.A0 (n_940) );
   OAI21X1 i_633 ( .Y (n_1035),
	.B0 (n_942),
	.A1 (n_911),
	.A0 (n_941) );
   OAI21X1 i_634 ( .Y (n_1036),
	.B0 (n_943),
	.A1 (n_912),
	.A0 (n_942) );
   OAI21X1 i_635 ( .Y (n_1037),
	.B0 (n_944),
	.A1 (n_913),
	.A0 (n_943) );
   OAI21X1 i_636 ( .Y (n_1038),
	.B0 (n_945),
	.A1 (n_914),
	.A0 (n_944) );
   OAI21X1 i_637 ( .Y (n_1039),
	.B0 (n_946),
	.A1 (n_915),
	.A0 (n_945) );
   OAI21X1 i_638 ( .Y (n_1040),
	.B0 (n_947),
	.A1 (n_916),
	.A0 (n_946) );
   OAI21X1 i_639 ( .Y (n_1041),
	.B0 (n_948),
	.A1 (n_917),
	.A0 (n_947) );
   OAI21X1 i_640 ( .Y (n_1042),
	.B0 (n_949),
	.A1 (n_918),
	.A0 (n_948) );
   OAI21X1 i_641 ( .Y (n_1043),
	.B0 (n_950),
	.A1 (n_919),
	.A0 (n_949) );
   OAI21X1 i_642 ( .Y (n_1044),
	.B0 (n_951),
	.A1 (n_920),
	.A0 (n_950) );
   OAI21X1 i_643 ( .Y (n_1045),
	.B0 (n_952),
	.A1 (n_921),
	.A0 (n_951) );
   OAI21X1 i_644 ( .Y (n_1046),
	.B0 (n_953),
	.A1 (n_922),
	.A0 (n_952) );
   OAI21X1 i_645 ( .Y (n_1047),
	.B0 (n_954),
	.A1 (n_923),
	.A0 (n_953) );
   OAI21X1 i_646 ( .Y (n_1048),
	.B0 (n_955),
	.A1 (n_924),
	.A0 (n_954) );
   OAI21X1 i_647 ( .Y (n_1049),
	.B0 (n_956),
	.A1 (n_925),
	.A0 (n_955) );
   OAI21X1 i_648 ( .Y (n_1050),
	.B0 (n_957),
	.A1 (n_926),
	.A0 (n_956) );
   OAI21X1 i_649 ( .Y (n_1051),
	.B0 (n_958),
	.A1 (n_927),
	.A0 (n_957) );
   OAI21X1 i_650 ( .Y (n_1052),
	.B0 (n_959),
	.A1 (n_928),
	.A0 (n_958) );
   OAI21X1 i_651 ( .Y (n_1053),
	.B0 (n_960),
	.A1 (n_929),
	.A0 (n_959) );
   AOI21X1 i_684 ( .Y (n_1086),
	.B0 (n_1026),
	.A1 (n_1056),
	.A0 (n_1024) );
   AOI21X1 i_685 ( .Y (n_1087),
	.B0 (n_1027),
	.A1 (n_1057),
	.A0 (n_1025) );
   AOI21X1 i_686 ( .Y (n_1088),
	.B0 (n_1028),
	.A1 (n_1058),
	.A0 (n_1026) );
   AOI21X1 i_687 ( .Y (n_1089),
	.B0 (n_1029),
	.A1 (n_1059),
	.A0 (n_1027) );
   AOI21X1 i_688 ( .Y (n_1090),
	.B0 (n_1030),
	.A1 (n_1060),
	.A0 (n_1028) );
   AOI21X1 i_689 ( .Y (n_1091),
	.B0 (n_1031),
	.A1 (n_1061),
	.A0 (n_1029) );
   AOI21X1 i_690 ( .Y (n_1092),
	.B0 (n_1032),
	.A1 (n_1062),
	.A0 (n_1030) );
   AOI21X1 i_691 ( .Y (n_1093),
	.B0 (n_1033),
	.A1 (n_1063),
	.A0 (n_1031) );
   AOI21X1 i_692 ( .Y (n_1094),
	.B0 (n_1034),
	.A1 (n_1064),
	.A0 (n_1032) );
   AOI21X1 i_693 ( .Y (n_1095),
	.B0 (n_1035),
	.A1 (n_1065),
	.A0 (n_1033) );
   AOI21X1 i_694 ( .Y (n_1096),
	.B0 (n_1036),
	.A1 (n_1066),
	.A0 (n_1034) );
   AOI21X1 i_695 ( .Y (n_1097),
	.B0 (n_1037),
	.A1 (n_1067),
	.A0 (n_1035) );
   AOI21X1 i_696 ( .Y (n_1098),
	.B0 (n_1038),
	.A1 (n_1068),
	.A0 (n_1036) );
   AOI21X1 i_697 ( .Y (n_1099),
	.B0 (n_1039),
	.A1 (n_1069),
	.A0 (n_1037) );
   AOI21X1 i_698 ( .Y (n_1100),
	.B0 (n_1040),
	.A1 (n_1070),
	.A0 (n_1038) );
   AOI21X1 i_699 ( .Y (n_1101),
	.B0 (n_1041),
	.A1 (n_1071),
	.A0 (n_1039) );
   AOI21X1 i_700 ( .Y (n_1102),
	.B0 (n_1042),
	.A1 (n_1072),
	.A0 (n_1040) );
   AOI21X1 i_701 ( .Y (n_1103),
	.B0 (n_1043),
	.A1 (n_1073),
	.A0 (n_1041) );
   AOI21X1 i_702 ( .Y (n_1104),
	.B0 (n_1044),
	.A1 (n_1074),
	.A0 (n_1042) );
   AOI21X1 i_703 ( .Y (n_1105),
	.B0 (n_1045),
	.A1 (n_1075),
	.A0 (n_1043) );
   AOI21X1 i_704 ( .Y (n_1106),
	.B0 (n_1046),
	.A1 (n_1076),
	.A0 (n_1044) );
   AOI21X1 i_705 ( .Y (n_1107),
	.B0 (n_1047),
	.A1 (n_1077),
	.A0 (n_1045) );
   AOI21X1 i_706 ( .Y (n_1108),
	.B0 (n_1048),
	.A1 (n_1078),
	.A0 (n_1046) );
   AOI21X1 i_707 ( .Y (n_1109),
	.B0 (n_1049),
	.A1 (n_1079),
	.A0 (n_1047) );
   AOI21X1 i_708 ( .Y (n_1110),
	.B0 (n_1050),
	.A1 (n_1080),
	.A0 (n_1048) );
   AOI21X1 i_709 ( .Y (n_1111),
	.B0 (n_1051),
	.A1 (n_1081),
	.A0 (n_1049) );
   AOI21X1 i_710 ( .Y (n_1112),
	.B0 (n_1052),
	.A1 (n_1082),
	.A0 (n_1050) );
   AOI21X1 i_711 ( .Y (n_1113),
	.B0 (n_1053),
	.A1 (n_1083),
	.A0 (n_1051) );
   OAI21X1 i_746 ( .Y (n_1148),
	.B0 (n_1088),
	.A1 (n_1118),
	.A0 (n_931) );
   OAI21X1 i_747 ( .Y (n_1149),
	.B0 (n_1089),
	.A1 (n_1119),
	.A0 (n_1085) );
   OAI21X1 i_748 ( .Y (n_1150),
	.B0 (n_1090),
	.A1 (n_1120),
	.A0 (n_1086) );
   OAI21X1 i_749 ( .Y (n_1151),
	.B0 (n_1091),
	.A1 (n_1121),
	.A0 (n_1087) );
   OAI21X1 i_750 ( .Y (n_1152),
	.B0 (n_1092),
	.A1 (n_1122),
	.A0 (n_1088) );
   OAI21X1 i_751 ( .Y (n_1153),
	.B0 (n_1093),
	.A1 (n_1123),
	.A0 (n_1089) );
   OAI21X1 i_752 ( .Y (n_1154),
	.B0 (n_1094),
	.A1 (n_1124),
	.A0 (n_1090) );
   OAI21X1 i_753 ( .Y (n_1155),
	.B0 (n_1095),
	.A1 (n_1125),
	.A0 (n_1091) );
   OAI21X1 i_754 ( .Y (n_1156),
	.B0 (n_1096),
	.A1 (n_1126),
	.A0 (n_1092) );
   OAI21X1 i_755 ( .Y (n_1157),
	.B0 (n_1097),
	.A1 (n_1127),
	.A0 (n_1093) );
   OAI21X1 i_756 ( .Y (n_1158),
	.B0 (n_1098),
	.A1 (n_1128),
	.A0 (n_1094) );
   OAI21X1 i_757 ( .Y (n_1159),
	.B0 (n_1099),
	.A1 (n_1129),
	.A0 (n_1095) );
   OAI21X1 i_758 ( .Y (n_1160),
	.B0 (n_1100),
	.A1 (n_1130),
	.A0 (n_1096) );
   OAI21X1 i_759 ( .Y (n_1161),
	.B0 (n_1101),
	.A1 (n_1131),
	.A0 (n_1097) );
   OAI21X1 i_760 ( .Y (n_1162),
	.B0 (n_1102),
	.A1 (n_1132),
	.A0 (n_1098) );
   OAI21X1 i_761 ( .Y (n_1163),
	.B0 (n_1103),
	.A1 (n_1133),
	.A0 (n_1099) );
   OAI21X1 i_762 ( .Y (n_1164),
	.B0 (n_1104),
	.A1 (n_1134),
	.A0 (n_1100) );
   OAI21X1 i_763 ( .Y (n_1165),
	.B0 (n_1105),
	.A1 (n_1135),
	.A0 (n_1101) );
   OAI21X1 i_764 ( .Y (n_1166),
	.B0 (n_1106),
	.A1 (n_1136),
	.A0 (n_1102) );
   OAI21X1 i_765 ( .Y (n_1167),
	.B0 (n_1107),
	.A1 (n_1137),
	.A0 (n_1103) );
   OAI21X1 i_766 ( .Y (n_1168),
	.B0 (n_1108),
	.A1 (n_1138),
	.A0 (n_1104) );
   OAI21X1 i_767 ( .Y (n_1169),
	.B0 (n_1109),
	.A1 (n_1139),
	.A0 (n_1105) );
   OAI21X1 i_768 ( .Y (n_1170),
	.B0 (n_1110),
	.A1 (n_1140),
	.A0 (n_1106) );
   OAI21X1 i_769 ( .Y (n_1171),
	.B0 (n_1111),
	.A1 (n_1141),
	.A0 (n_1107) );
   OAI21X1 i_770 ( .Y (n_1172),
	.B0 (n_1112),
	.A1 (n_1142),
	.A0 (n_1108) );
   OAI21X1 i_771 ( .Y (n_1173),
	.B0 (n_1113),
	.A1 (n_1143),
	.A0 (n_1109) );
   AOI21X1 i_810 ( .Y (n_1212),
	.B0 (n_1152),
	.A1 (n_1182),
	.A0 (n_1024) );
   AOI21X1 i_811 ( .Y (n_1213),
	.B0 (n_1153),
	.A1 (n_1183),
	.A0 (n_1025) );
   AOI21X1 i_812 ( .Y (n_1214),
	.B0 (n_1154),
	.A1 (n_1184),
	.A0 (n_1146) );
   AOI21X1 i_813 ( .Y (n_1215),
	.B0 (n_1155),
	.A1 (n_1185),
	.A0 (n_1147) );
   AOI21X1 i_814 ( .Y (n_1216),
	.B0 (n_1156),
	.A1 (n_1186),
	.A0 (n_1148) );
   AOI21X1 i_815 ( .Y (n_1217),
	.B0 (n_1157),
	.A1 (n_1187),
	.A0 (n_1149) );
   AOI21X1 i_816 ( .Y (n_1218),
	.B0 (n_1158),
	.A1 (n_1188),
	.A0 (n_1150) );
   AOI21X1 i_817 ( .Y (n_1219),
	.B0 (n_1159),
	.A1 (n_1189),
	.A0 (n_1151) );
   AOI21X1 i_818 ( .Y (n_1220),
	.B0 (n_1160),
	.A1 (n_1190),
	.A0 (n_1152) );
   AOI21X1 i_819 ( .Y (n_1221),
	.B0 (n_1161),
	.A1 (n_1191),
	.A0 (n_1153) );
   AOI21X1 i_820 ( .Y (n_1222),
	.B0 (n_1162),
	.A1 (n_1192),
	.A0 (n_1154) );
   AOI21X1 i_821 ( .Y (n_1223),
	.B0 (n_1163),
	.A1 (n_1193),
	.A0 (n_1155) );
   AOI21X1 i_822 ( .Y (n_1224),
	.B0 (n_1164),
	.A1 (n_1194),
	.A0 (n_1156) );
   AOI21X1 i_823 ( .Y (n_1225),
	.B0 (n_1165),
	.A1 (n_1195),
	.A0 (n_1157) );
   AOI21X1 i_824 ( .Y (n_1226),
	.B0 (n_1166),
	.A1 (n_1196),
	.A0 (n_1158) );
   AOI21X1 i_825 ( .Y (n_1227),
	.B0 (n_1167),
	.A1 (n_1197),
	.A0 (n_1159) );
   AOI21X1 i_826 ( .Y (n_1228),
	.B0 (n_1168),
	.A1 (n_1198),
	.A0 (n_1160) );
   AOI21X1 i_827 ( .Y (n_1229),
	.B0 (n_1169),
	.A1 (n_1199),
	.A0 (n_1161) );
   AOI21X1 i_828 ( .Y (n_1230),
	.B0 (n_1170),
	.A1 (n_1200),
	.A0 (n_1162) );
   AOI21X1 i_829 ( .Y (n_1231),
	.B0 (n_1171),
	.A1 (n_1201),
	.A0 (n_1163) );
   AOI21X1 i_830 ( .Y (n_1232),
	.B0 (n_1172),
	.A1 (n_1202),
	.A0 (n_1164) );
   AOI21X1 i_831 ( .Y (n_1233),
	.B0 (n_1173),
	.A1 (n_1203),
	.A0 (n_1165) );
   OAI21X1 i_878 ( .Y (n_1280),
	.B0 (n_1220),
	.A1 (n_1250),
	.A0 (n_931) );
   OAI21X1 i_879 ( .Y (n_1281),
	.B0 (n_1221),
	.A1 (n_1251),
	.A0 (n_1085) );
   OAI21X1 i_880 ( .Y (n_1282),
	.B0 (n_1222),
	.A1 (n_1252),
	.A0 (n_1086) );
   OAI21X1 i_881 ( .Y (n_1283),
	.B0 (n_1223),
	.A1 (n_1253),
	.A0 (n_1087) );
   OAI21X1 i_882 ( .Y (n_1284),
	.B0 (n_1224),
	.A1 (n_1254),
	.A0 (n_1208) );
   OAI21X1 i_883 ( .Y (n_1285),
	.B0 (n_1225),
	.A1 (n_1255),
	.A0 (n_1209) );
   OAI21X1 i_884 ( .Y (n_1286),
	.B0 (n_1226),
	.A1 (n_1256),
	.A0 (n_1210) );
   OAI21X1 i_885 ( .Y (n_1287),
	.B0 (n_1227),
	.A1 (n_1257),
	.A0 (n_1211) );
   OAI21X1 i_886 ( .Y (n_1288),
	.B0 (n_1228),
	.A1 (n_1258),
	.A0 (n_1212) );
   OAI21X1 i_887 ( .Y (n_1289),
	.B0 (n_1229),
	.A1 (n_1259),
	.A0 (n_1213) );
   OAI21X1 i_888 ( .Y (n_1290),
	.B0 (n_1230),
	.A1 (n_1260),
	.A0 (n_1214) );
   OAI21X1 i_889 ( .Y (n_1291),
	.B0 (n_1231),
	.A1 (n_1261),
	.A0 (n_1215) );
   OAI21X1 i_890 ( .Y (n_1292),
	.B0 (n_1232),
	.A1 (n_1262),
	.A0 (n_1216) );
   OAI21X1 i_891 ( .Y (y[31]),
	.B0 (n_1233),
	.A1 (n_1263),
	.A0 (n_1217) );
endmodule

module mult_32 (
	ovm,
	op_a,
	op_b,
	result );
   input ovm;
   input [15:0] op_a;
   input [15:0] op_b;
   output [31:0] result;

   // Internal wires
   wire \ab_result[22] ;
   wire n_588;
   wire n_361;
   wire \ab_result[23] ;
   wire n_587;
   wire n_359;
   wire \ab_result[24] ;
   wire n_586;
   wire \ab_result[25] ;
   wire n_3099;
   wire n_354;
   wire \ab_result[26] ;
   wire n_584;
   wire n_351;
   wire \ab_result[27] ;
   wire n_583;
   wire n_348;
   wire \ab_result[28] ;
   wire n_582;
   wire n_345;
   wire n_579;
   wire n_520;
   wire n_545;
   wire n_577;
   wire n_344;
   wire \ab_result[29] ;
   wire n_564;
   wire \ab_result[30] ;
   wire n_549;
   wire \ab_result[31] ;
   wire n_527;
   wire n_336;
   wire n_334;
   wire n_333;
   wire n_497;
   wire n_331;
   wire \ab_b[1] ;
   wire n_496;
   wire n_329;
   wire \ab_b[2] ;
   wire n_495;
   wire n_327;
   wire \ab_b[3] ;
   wire n_494;
   wire n_325;
   wire \ab_b[4] ;
   wire n_493;
   wire n_322;
   wire \ab_b[5] ;
   wire n_492;
   wire n_320;
   wire \ab_b[6] ;
   wire n_491;
   wire n_318;
   wire \ab_b[7] ;
   wire n_490;
   wire n_316;
   wire \ab_b[8] ;
   wire n_489;
   wire n_314;
   wire \ab_b[9] ;
   wire n_488;
   wire n_312;
   wire \ab_b[10] ;
   wire n_487;
   wire n_310;
   wire \ab_b[11] ;
   wire n_486;
   wire n_308;
   wire \ab_b[12] ;
   wire n_479;
   wire n_305;
   wire \ab_b[13] ;
   wire n_474;
   wire n_302;
   wire \ab_b[14] ;
   wire n_451;
   wire n_299;
   wire \ab_a[1] ;
   wire n_450;
   wire n_297;
   wire \ab_a[2] ;
   wire n_449;
   wire n_295;
   wire \ab_a[3] ;
   wire n_448;
   wire n_293;
   wire \ab_a[4] ;
   wire n_447;
   wire n_290;
   wire \ab_a[5] ;
   wire n_446;
   wire n_288;
   wire \ab_a[6] ;
   wire n_445;
   wire n_286;
   wire \ab_a[7] ;
   wire n_444;
   wire n_284;
   wire \ab_a[8] ;
   wire n_443;
   wire n_282;
   wire \ab_a[9] ;
   wire n_442;
   wire n_280;
   wire \ab_a[10] ;
   wire n_441;
   wire n_278;
   wire \ab_a[11] ;
   wire n_440;
   wire n_276;
   wire \ab_a[12] ;
   wire n_433;
   wire n_273;
   wire \ab_a[13] ;
   wire n_428;
   wire n_270;
   wire \ab_a[14] ;
   wire n_268;
   wire n_558;
   wire \ab_result[21] ;
   wire n_363;
   wire \ab_result[20] ;
   wire n_365;
   wire n_515;
   wire \ab_result[19] ;
   wire n_367;
   wire n_539;
   wire \ab_result[18] ;
   wire n_369;
   wire \ab_result[17] ;
   wire n_593;
   wire \ab_result[16] ;
   wire n_594;
   wire \ab_result[15] ;
   wire n_595;
   wire \ab_result[14] ;
   wire n_596;
   wire n_554;
   wire \ab_result[13] ;
   wire n_379;
   wire n_571;
   wire \ab_result[12] ;
   wire n_381;
   wire n_507;
   wire \ab_result[11] ;
   wire n_383;
   wire n_533;
   wire \ab_result[10] ;
   wire n_385;
   wire \ab_result[9] ;
   wire n_601;
   wire n_387;
   wire \ab_result[8] ;
   wire n_602;
   wire \ab_result[7] ;
   wire n_603;
   wire \ab_result[6] ;
   wire n_604;
   wire \ab_result[5] ;
   wire n_605;
   wire n_499;
   wire \ab_result[3] ;
   wire n_397;
   wire \ab_result[4] ;
   wire n_398;
   wire n_400;
   wire n_498;
   wire \ab_result[2] ;
   wire n_402;
   wire \ab_result[1] ;
   wire n_609;
   wire n_404;
   wire n_406;
   wire n_407;
   wire n_408;
   wire n_409;
   wire n_3101;
   wire n_411;
   wire n_412;
   wire n_413;
   wire n_415;
   wire n_416;
   wire n_417;
   wire n_420;
   wire n_422;
   wire n_425;
   wire n_427;
   wire n_429;
   wire n_431;
   wire n_432;
   wire n_435;
   wire n_437;
   wire n_439;
   wire n_452;
   wire n_453;
   wire n_454;
   wire n_455;
   wire n_3100;
   wire n_457;
   wire n_458;
   wire n_459;
   wire n_461;
   wire n_462;
   wire n_463;
   wire n_466;
   wire n_468;
   wire n_471;
   wire n_473;
   wire n_475;
   wire n_477;
   wire n_478;
   wire n_481;
   wire n_483;
   wire n_485;
   wire n_500;
   wire n_501;
   wire n_503;
   wire n_504;
   wire n_505;
   wire n_508;
   wire n_509;
   wire n_511;
   wire n_512;
   wire n_513;
   wire n_516;
   wire n_517;
   wire n_519;
   wire n_522;
   wire n_525;
   wire n_528;
   wire n_530;
   wire n_534;
   wire n_536;
   wire n_541;
   wire n_542;
   wire n_544;
   wire n_548;
   wire n_552;
   wire n_556;
   wire n_560;
   wire n_562;
   wire n_566;
   wire n_568;
   wire n_572;
   wire n_574;
   wire n_578;
   wire n_585;
   wire \ab_a[15] ;
   wire \ab_b[15] ;

   OAI21XL i_818589 ( .Y (result[22]),
	.B0 (n_361),
	.A1 (n_588),
	.A0 (\ab_result[22] ) );
   NAND2X1 i_320 ( .Y (n_361),
	.B (n_588),
	.A (\ab_result[22] ) );
   OAI21XL i_808588 ( .Y (result[23]),
	.B0 (n_359),
	.A1 (n_587),
	.A0 (\ab_result[23] ) );
   NAND2X1 i_317 ( .Y (n_359),
	.B (n_587),
	.A (\ab_result[23] ) );
   XOR2X1 i_798587 ( .Y (result[24]),
	.B (n_586),
	.A (\ab_result[24] ) );
   OAI21XL i_788586 ( .Y (result[25]),
	.B0 (n_354),
	.A1 (n_3099),
	.A0 (\ab_result[25] ) );
   NAND2X1 i_310 ( .Y (n_354),
	.B (n_3099),
	.A (\ab_result[25] ) );
   OAI21XL i_778585 ( .Y (result[26]),
	.B0 (n_351),
	.A1 (n_584),
	.A0 (\ab_result[26] ) );
   NAND2X1 i_306 ( .Y (n_351),
	.B (n_584),
	.A (\ab_result[26] ) );
   OAI21XL i_768584 ( .Y (result[27]),
	.B0 (n_348),
	.A1 (n_583),
	.A0 (\ab_result[27] ) );
   NAND2X1 i_302 ( .Y (n_348),
	.B (n_583),
	.A (\ab_result[27] ) );
   OAI21XL i_758583 ( .Y (result[28]),
	.B0 (n_345),
	.A1 (n_582),
	.A0 (\ab_result[28] ) );
   NAND2X1 i_298 ( .Y (n_345),
	.B (n_582),
	.A (\ab_result[28] ) );
   NAND4BXL i_295 ( .Y (n_344),
	.D (n_577),
	.C (n_545),
	.B (n_520),
	.AN (n_579) );
   XOR2X1 i_748582 ( .Y (result[29]),
	.B (n_564),
	.A (\ab_result[29] ) );
   XOR2X1 i_738581 ( .Y (result[30]),
	.B (n_549),
	.A (\ab_result[30] ) );
   OAI21XL i_728580 ( .Y (result[31]),
	.B0 (n_336),
	.A1 (n_527),
	.A0 (\ab_result[31] ) );
   NAND2X1 i_250 ( .Y (n_336),
	.B (n_527),
	.A (\ab_result[31] ) );
   NOR2BX1 i_238 ( .Y (n_334),
	.B (op_b[15]),
	.AN (op_a[15]) );
   NOR2BX1 i_237 ( .Y (n_333),
	.B (op_a[15]),
	.AN (op_b[15]) );
   OAI21XL i_388412 ( .Y (\ab_b[1] ),
	.B0 (n_331),
	.A1 (n_497),
	.A0 (op_b[1]) );
   NAND2X1 i_234 ( .Y (n_331),
	.B (n_497),
	.A (op_b[1]) );
   OAI21XL i_378411 ( .Y (\ab_b[2] ),
	.B0 (n_329),
	.A1 (n_496),
	.A0 (op_b[2]) );
   NAND2X1 i_231 ( .Y (n_329),
	.B (n_496),
	.A (op_b[2]) );
   OAI21XL i_368410 ( .Y (\ab_b[3] ),
	.B0 (n_327),
	.A1 (n_495),
	.A0 (op_b[3]) );
   NAND2X1 i_228 ( .Y (n_327),
	.B (n_495),
	.A (op_b[3]) );
   OAI21XL i_358409 ( .Y (\ab_b[4] ),
	.B0 (n_325),
	.A1 (n_494),
	.A0 (op_b[4]) );
   NAND2X1 i_225 ( .Y (n_325),
	.B (n_494),
	.A (op_b[4]) );
   OAI21XL i_348408 ( .Y (\ab_b[5] ),
	.B0 (n_322),
	.A1 (n_493),
	.A0 (op_b[5]) );
   NAND2X1 i_221 ( .Y (n_322),
	.B (n_493),
	.A (op_b[5]) );
   OAI21XL i_338407 ( .Y (\ab_b[6] ),
	.B0 (n_320),
	.A1 (n_492),
	.A0 (op_b[6]) );
   NAND2X1 i_218 ( .Y (n_320),
	.B (n_492),
	.A (op_b[6]) );
   OAI21XL i_328406 ( .Y (\ab_b[7] ),
	.B0 (n_318),
	.A1 (n_491),
	.A0 (op_b[7]) );
   NAND2X1 i_215 ( .Y (n_318),
	.B (n_491),
	.A (op_b[7]) );
   OAI21XL i_318405 ( .Y (\ab_b[8] ),
	.B0 (n_316),
	.A1 (n_490),
	.A0 (op_b[8]) );
   NAND2X1 i_212 ( .Y (n_316),
	.B (n_490),
	.A (op_b[8]) );
   OAI21XL i_308404 ( .Y (\ab_b[9] ),
	.B0 (n_314),
	.A1 (n_489),
	.A0 (op_b[9]) );
   NAND2X1 i_209 ( .Y (n_314),
	.B (n_489),
	.A (op_b[9]) );
   OAI21XL i_298403 ( .Y (\ab_b[10] ),
	.B0 (n_312),
	.A1 (n_488),
	.A0 (op_b[10]) );
   NAND2X1 i_206 ( .Y (n_312),
	.B (n_488),
	.A (op_b[10]) );
   OAI21XL i_288402 ( .Y (\ab_b[11] ),
	.B0 (n_310),
	.A1 (n_487),
	.A0 (op_b[11]) );
   NAND2X1 i_203 ( .Y (n_310),
	.B (n_487),
	.A (op_b[11]) );
   OAI21XL i_278401 ( .Y (\ab_b[12] ),
	.B0 (n_308),
	.A1 (n_486),
	.A0 (op_b[12]) );
   NAND2X1 i_200 ( .Y (n_308),
	.B (n_486),
	.A (op_b[12]) );
   OAI21XL i_268400 ( .Y (\ab_b[13] ),
	.B0 (n_305),
	.A1 (n_479),
	.A0 (op_b[13]) );
   NAND2X1 i_191 ( .Y (n_305),
	.B (n_479),
	.A (op_b[13]) );
   OAI21XL i_258399 ( .Y (\ab_b[14] ),
	.B0 (n_302),
	.A1 (n_474),
	.A0 (op_b[14]) );
   NAND2X1 i_183 ( .Y (n_302),
	.B (n_474),
	.A (op_b[14]) );
   OAI21XL i_388364 ( .Y (\ab_a[1] ),
	.B0 (n_299),
	.A1 (n_451),
	.A0 (op_a[1]) );
   NAND2X1 i_168 ( .Y (n_299),
	.B (n_451),
	.A (op_a[1]) );
   OAI21XL i_378363 ( .Y (\ab_a[2] ),
	.B0 (n_297),
	.A1 (n_450),
	.A0 (op_a[2]) );
   NAND2X1 i_165 ( .Y (n_297),
	.B (n_450),
	.A (op_a[2]) );
   OAI21XL i_368362 ( .Y (\ab_a[3] ),
	.B0 (n_295),
	.A1 (n_449),
	.A0 (op_a[3]) );
   NAND2X1 i_162 ( .Y (n_295),
	.B (n_449),
	.A (op_a[3]) );
   OAI21XL i_358361 ( .Y (\ab_a[4] ),
	.B0 (n_293),
	.A1 (n_448),
	.A0 (op_a[4]) );
   NAND2X1 i_159 ( .Y (n_293),
	.B (n_448),
	.A (op_a[4]) );
   OAI21XL i_348360 ( .Y (\ab_a[5] ),
	.B0 (n_290),
	.A1 (n_447),
	.A0 (op_a[5]) );
   NAND2X1 i_155 ( .Y (n_290),
	.B (n_447),
	.A (op_a[5]) );
   OAI21XL i_338359 ( .Y (\ab_a[6] ),
	.B0 (n_288),
	.A1 (n_446),
	.A0 (op_a[6]) );
   NAND2X1 i_152 ( .Y (n_288),
	.B (n_446),
	.A (op_a[6]) );
   OAI21XL i_328358 ( .Y (\ab_a[7] ),
	.B0 (n_286),
	.A1 (n_445),
	.A0 (op_a[7]) );
   NAND2X1 i_142 ( .Y (n_286),
	.B (n_445),
	.A (op_a[7]) );
   OAI21XL i_318357 ( .Y (\ab_a[8] ),
	.B0 (n_284),
	.A1 (n_444),
	.A0 (op_a[8]) );
   NAND2X1 i_139 ( .Y (n_284),
	.B (n_444),
	.A (op_a[8]) );
   OAI21XL i_308356 ( .Y (\ab_a[9] ),
	.B0 (n_282),
	.A1 (n_443),
	.A0 (op_a[9]) );
   NAND2X1 i_136 ( .Y (n_282),
	.B (n_443),
	.A (op_a[9]) );
   OAI21XL i_298355 ( .Y (\ab_a[10] ),
	.B0 (n_280),
	.A1 (n_442),
	.A0 (op_a[10]) );
   NAND2X1 i_133 ( .Y (n_280),
	.B (n_442),
	.A (op_a[10]) );
   OAI21XL i_288354 ( .Y (\ab_a[11] ),
	.B0 (n_278),
	.A1 (n_441),
	.A0 (op_a[11]) );
   NAND2X1 i_130 ( .Y (n_278),
	.B (n_441),
	.A (op_a[11]) );
   OAI21XL i_278353 ( .Y (\ab_a[12] ),
	.B0 (n_276),
	.A1 (n_440),
	.A0 (op_a[12]) );
   NAND2X1 i_127 ( .Y (n_276),
	.B (n_440),
	.A (op_a[12]) );
   OAI21XL i_268352 ( .Y (\ab_a[13] ),
	.B0 (n_273),
	.A1 (n_433),
	.A0 (op_a[13]) );
   NAND2X1 i_118 ( .Y (n_273),
	.B (n_433),
	.A (op_a[13]) );
   OAI21XL i_258351 ( .Y (\ab_a[14] ),
	.B0 (n_270),
	.A1 (n_428),
	.A0 (op_a[14]) );
   NAND2X1 i_102 ( .Y (n_270),
	.B (n_428),
	.A (op_a[14]) );
   NOR2X1 i_6286 ( .Y (n_268),
	.B (n_333),
	.A (n_334) );
   OAI21XL i_323 ( .Y (n_363),
	.B0 (\ab_result[21] ),
	.A1 (n_268),
	.A0 (n_558) );
   OAI31X1 i_828590 ( .Y (result[21]),
	.B0 (n_363),
	.A2 (n_558),
	.A1 (\ab_result[21] ),
	.A0 (n_268) );
   OAI21XL i_326 ( .Y (n_365),
	.B0 (\ab_result[20] ),
	.A1 (n_268),
	.A0 (n_577) );
   OAI31X1 i_838591 ( .Y (result[20]),
	.B0 (n_365),
	.A2 (n_268),
	.A1 (\ab_result[20] ),
	.A0 (n_577) );
   OAI21XL i_329 ( .Y (n_367),
	.B0 (\ab_result[19] ),
	.A1 (n_268),
	.A0 (n_515) );
   OAI31X1 i_848592 ( .Y (result[19]),
	.B0 (n_367),
	.A2 (n_515),
	.A1 (\ab_result[19] ),
	.A0 (n_268) );
   OAI21XL i_332 ( .Y (n_369),
	.B0 (\ab_result[18] ),
	.A1 (n_268),
	.A0 (n_539) );
   OAI31X1 i_858593 ( .Y (result[18]),
	.B0 (n_369),
	.A2 (\ab_result[18] ),
	.A1 (n_268),
	.A0 (n_539) );
   XOR2X1 i_868594 ( .Y (result[17]),
	.B (n_593),
	.A (\ab_result[17] ) );
   XOR2X1 i_878595 ( .Y (result[16]),
	.B (n_594),
	.A (\ab_result[16] ) );
   XOR2X1 i_888596 ( .Y (result[15]),
	.B (n_595),
	.A (\ab_result[15] ) );
   XOR2X1 i_898597 ( .Y (result[14]),
	.B (n_596),
	.A (\ab_result[14] ) );
   OAI21XL i_347 ( .Y (n_379),
	.B0 (\ab_result[13] ),
	.A1 (n_268),
	.A0 (n_554) );
   OAI31X1 i_908598 ( .Y (result[13]),
	.B0 (n_379),
	.A2 (n_554),
	.A1 (\ab_result[13] ),
	.A0 (n_268) );
   OAI21XL i_350 ( .Y (n_381),
	.B0 (\ab_result[12] ),
	.A1 (n_268),
	.A0 (n_571) );
   OAI31X1 i_918599 ( .Y (result[12]),
	.B0 (n_381),
	.A2 (\ab_result[12] ),
	.A1 (n_268),
	.A0 (n_571) );
   OAI21XL i_353 ( .Y (n_383),
	.B0 (\ab_result[11] ),
	.A1 (n_268),
	.A0 (n_507) );
   OAI31X1 i_928600 ( .Y (result[11]),
	.B0 (n_383),
	.A2 (n_507),
	.A1 (\ab_result[11] ),
	.A0 (n_268) );
   OAI21XL i_356 ( .Y (n_385),
	.B0 (\ab_result[10] ),
	.A1 (n_268),
	.A0 (n_533) );
   OAI31X1 i_938601 ( .Y (result[10]),
	.B0 (n_385),
	.A2 (\ab_result[10] ),
	.A1 (n_268),
	.A0 (n_533) );
   NAND2X1 i_359 ( .Y (n_387),
	.B (n_601),
	.A (\ab_result[9] ) );
   OAI21XL i_948602 ( .Y (result[9]),
	.B0 (n_387),
	.A1 (n_601),
	.A0 (\ab_result[9] ) );
   XOR2X1 i_95 ( .Y (result[8]),
	.B (n_602),
	.A (\ab_result[8] ) );
   XOR2X1 i_968603 ( .Y (result[7]),
	.B (n_603),
	.A (\ab_result[7] ) );
   XOR2X1 i_97 ( .Y (result[6]),
	.B (n_604),
	.A (\ab_result[6] ) );
   XOR2X1 i_98 ( .Y (result[5]),
	.B (n_605),
	.A (\ab_result[5] ) );
   NOR2BX1 i_374 ( .Y (n_397),
	.B (\ab_result[3] ),
	.AN (n_499) );
   OAI21XL i_375 ( .Y (n_398),
	.B0 (\ab_result[4] ),
	.A1 (n_268),
	.A0 (n_397) );
   OAI31X1 i_998604 ( .Y (result[4]),
	.B0 (n_398),
	.A2 (n_397),
	.A1 (\ab_result[4] ),
	.A0 (n_268) );
   OAI21XL i_378 ( .Y (n_400),
	.B0 (\ab_result[3] ),
	.A1 (n_268),
	.A0 (n_499) );
   OAI31X1 i_1008605 ( .Y (result[3]),
	.B0 (n_400),
	.A2 (\ab_result[3] ),
	.A1 (n_268),
	.A0 (n_499) );
   OAI21XL i_381 ( .Y (n_402),
	.B0 (\ab_result[2] ),
	.A1 (n_268),
	.A0 (n_498) );
   OAI31X1 i_1018606 ( .Y (result[2]),
	.B0 (n_402),
	.A2 (\ab_result[2] ),
	.A1 (n_268),
	.A0 (n_498) );
   NAND2X1 i_384 ( .Y (n_404),
	.B (n_609),
	.A (\ab_result[1] ) );
   OAI21XL i_1028607 ( .Y (result[1]),
	.B0 (n_404),
	.A1 (n_609),
	.A0 (\ab_result[1] ) );
   NOR2X1 i_1 ( .Y (n_406),
	.B (op_a[0]),
	.A (op_a[1]) );
   NAND2BX1 i_181705 ( .Y (n_407),
	.B (n_406),
	.AN (op_a[2]) );
   NOR2X1 i_39 ( .Y (n_408),
	.B (op_a[4]),
	.A (op_a[3]) );
   NOR2X1 i_40 ( .Y (n_409),
	.B (op_a[6]),
	.A (op_a[5]) );
   NAND3X1 i_381723 ( .Y (n_411),
	.C (n_3101),
	.B (n_409),
	.A (n_408) );
   NOR2X1 i_25 ( .Y (n_412),
	.B (op_a[8]),
	.A (op_a[7]) );
   NOR2X1 i_41 ( .Y (n_413),
	.B (op_a[10]),
	.A (op_a[9]) );
   NOR4BX1 i_58 ( .Y (n_415),
	.D (n_411),
	.C (op_a[8]),
	.B (op_a[7]),
	.AN (n_413) );
   NOR2X1 i_24 ( .Y (n_416),
	.B (op_a[12]),
	.A (op_a[11]) );
   NOR2X1 i_89 ( .Y (n_417),
	.B (op_a[14]),
	.A (op_a[13]) );
   NOR2X1 i_92 ( .Y (n_420),
	.B (op_a[5]),
	.A (op_a[2]) );
   NAND3X1 i_371722 ( .Y (n_422),
	.C (n_406),
	.B (n_420),
	.A (n_408) );
   NOR4BX1 i_57 ( .Y (n_425),
	.D (n_422),
	.C (op_a[9]),
	.B (op_a[6]),
	.AN (n_412) );
   NOR4X1 i_101 ( .Y (n_427),
	.D (op_a[13]),
	.C (op_a[10]),
	.B (op_a[12]),
	.A (op_a[11]) );
   OAI2BB1X1 i_3 ( .Y (n_428),
	.B0 (op_a[15]),
	.A1N (n_427),
	.A0N (n_425) );
   NAND2X1 i_361721 ( .Y (n_429),
	.B (n_3101),
	.A (n_408) );
   NAND4X1 i_56 ( .Y (n_431),
	.D (n_3101),
	.C (n_412),
	.B (n_409),
	.A (n_408) );
   NAND2X1 i_117 ( .Y (n_432),
	.B (n_416),
	.A (n_413) );
   OAI21XL i_4 ( .Y (n_433),
	.B0 (op_a[15]),
	.A1 (n_432),
	.A0 (n_431) );
   NOR3X1 i_122 ( .Y (n_435),
	.C (op_a[3]),
	.B (op_a[7]),
	.A (op_a[4]) );
   NAND3X1 i_09003 ( .Y (n_437),
	.C (n_3101),
	.B (n_435),
	.A (n_409) );
   OR4X1 i_126 ( .Y (n_439),
	.D (op_a[11]),
	.C (op_a[8]),
	.B (op_a[10]),
	.A (op_a[9]) );
   OAI21XL i_5 ( .Y (n_440),
	.B0 (op_a[15]),
	.A1 (n_439),
	.A0 (n_437) );
   NAND2BX1 i_42 ( .Y (n_441),
	.B (op_a[15]),
	.AN (n_415) );
   NAND2BX1 i_43 ( .Y (n_442),
	.B (op_a[15]),
	.AN (n_425) );
   NAND2X1 i_44 ( .Y (n_443),
	.B (n_431),
	.A (op_a[15]) );
   NAND2X1 i_45 ( .Y (n_444),
	.B (n_437),
	.A (op_a[15]) );
   NAND2X1 i_46 ( .Y (n_445),
	.B (n_411),
	.A (op_a[15]) );
   NAND2X1 i_47 ( .Y (n_446),
	.B (n_422),
	.A (op_a[15]) );
   NAND2X1 i_48 ( .Y (n_447),
	.B (n_429),
	.A (op_a[15]) );
   OAI21XL i_6 ( .Y (n_448),
	.B0 (op_a[15]),
	.A1 (n_407),
	.A0 (op_a[3]) );
   NAND2X1 i_49 ( .Y (n_449),
	.B (n_407),
	.A (op_a[15]) );
   OAI21XL i_50 ( .Y (n_450),
	.B0 (op_a[15]),
	.A1 (op_a[0]),
	.A0 (op_a[1]) );
   NAND2X1 i_51 ( .Y (n_451),
	.B (op_a[0]),
	.A (op_a[15]) );
   NOR2X1 i_11967 ( .Y (n_452),
	.B (op_b[0]),
	.A (op_b[1]) );
   NAND2BX1 i_181983 ( .Y (n_453),
	.B (n_452),
	.AN (op_b[2]) );
   NOR2X1 i_36 ( .Y (n_454),
	.B (op_b[4]),
	.A (op_b[3]) );
   NOR2X1 i_37 ( .Y (n_455),
	.B (op_b[6]),
	.A (op_b[5]) );
   NAND3X1 i_382001 ( .Y (n_457),
	.C (n_3100),
	.B (n_455),
	.A (n_454) );
   NOR2X1 i_22 ( .Y (n_458),
	.B (op_b[8]),
	.A (op_b[7]) );
   NOR2X1 i_38 ( .Y (n_459),
	.B (op_b[10]),
	.A (op_b[9]) );
   NOR4BX1 i_582018 ( .Y (n_461),
	.D (n_457),
	.C (op_b[8]),
	.B (op_b[7]),
	.AN (n_459) );
   NOR2X1 i_23 ( .Y (n_462),
	.B (op_b[12]),
	.A (op_b[11]) );
   NOR2X1 i_173 ( .Y (n_463),
	.B (op_b[14]),
	.A (op_b[13]) );
   NOR2X1 i_176 ( .Y (n_466),
	.B (op_b[5]),
	.A (op_b[2]) );
   NAND3X1 i_372000 ( .Y (n_468),
	.C (n_452),
	.B (n_466),
	.A (n_454) );
   NOR4BX1 i_572017 ( .Y (n_471),
	.D (n_468),
	.C (op_b[9]),
	.B (op_b[6]),
	.AN (n_458) );
   NOR4X1 i_182 ( .Y (n_473),
	.D (op_b[13]),
	.C (op_b[10]),
	.B (op_b[12]),
	.A (op_b[11]) );
   OAI2BB1X1 i_7 ( .Y (n_474),
	.B0 (op_b[15]),
	.A1N (n_473),
	.A0N (n_471) );
   NAND2X1 i_361999 ( .Y (n_475),
	.B (n_3100),
	.A (n_454) );
   NAND4X1 i_562016 ( .Y (n_477),
	.D (n_3100),
	.C (n_458),
	.B (n_455),
	.A (n_454) );
   NAND2X1 i_190 ( .Y (n_478),
	.B (n_462),
	.A (n_459) );
   OAI21XL i_8 ( .Y (n_479),
	.B0 (op_b[15]),
	.A1 (n_478),
	.A0 (n_477) );
   NOR3X1 i_195 ( .Y (n_481),
	.C (op_b[3]),
	.B (op_b[7]),
	.A (op_b[4]) );
   NAND3X1 i_2 ( .Y (n_483),
	.C (n_3100),
	.B (n_481),
	.A (n_455) );
   OR4X1 i_199 ( .Y (n_485),
	.D (op_b[11]),
	.C (op_b[8]),
	.B (op_b[10]),
	.A (op_b[9]) );
   OAI21XL i_9 ( .Y (n_486),
	.B0 (op_b[15]),
	.A1 (n_485),
	.A0 (n_483) );
   NAND2BX1 i_52 ( .Y (n_487),
	.B (op_b[15]),
	.AN (n_461) );
   NAND2BX1 i_53 ( .Y (n_488),
	.B (op_b[15]),
	.AN (n_471) );
   NAND2X1 i_54 ( .Y (n_489),
	.B (n_477),
	.A (op_b[15]) );
   NAND2X1 i_55 ( .Y (n_490),
	.B (n_483),
	.A (op_b[15]) );
   NAND2X1 i_59 ( .Y (n_491),
	.B (n_457),
	.A (op_b[15]) );
   NAND2X1 i_60 ( .Y (n_492),
	.B (n_468),
	.A (op_b[15]) );
   NAND2X1 i_61 ( .Y (n_493),
	.B (n_475),
	.A (op_b[15]) );
   OAI21XL i_10 ( .Y (n_494),
	.B0 (op_b[15]),
	.A1 (n_453),
	.A0 (op_b[3]) );
   NAND2X1 i_62 ( .Y (n_495),
	.B (n_453),
	.A (op_b[15]) );
   OAI21XL i_63 ( .Y (n_496),
	.B0 (op_b[15]),
	.A1 (op_b[0]),
	.A0 (op_b[1]) );
   NAND2X1 i_64 ( .Y (n_497),
	.B (op_b[0]),
	.A (op_b[15]) );
   NOR2X1 i_12117 ( .Y (n_498),
	.B (result[0]),
	.A (\ab_result[1] ) );
   NOR3X1 i_342149 ( .Y (n_499),
	.C (\ab_result[2] ),
	.B (result[0]),
	.A (\ab_result[1] ) );
   NOR2X1 i_26 ( .Y (n_500),
	.B (\ab_result[4] ),
	.A (\ab_result[3] ) );
   NOR2X1 i_27 ( .Y (n_501),
	.B (\ab_result[6] ),
	.A (\ab_result[5] ) );
   NAND3X1 i_702180 ( .Y (n_503),
	.C (n_499),
	.B (n_501),
	.A (n_500) );
   NOR2X1 i_28 ( .Y (n_504),
	.B (\ab_result[8] ),
	.A (\ab_result[7] ) );
   NOR2X1 i_29 ( .Y (n_505),
	.B (\ab_result[10] ),
	.A (\ab_result[9] ) );
   NOR4BX1 i_106 ( .Y (n_507),
	.D (n_503),
	.C (\ab_result[8] ),
	.B (\ab_result[7] ),
	.AN (n_505) );
   NOR2X1 i_30 ( .Y (n_508),
	.B (\ab_result[12] ),
	.A (\ab_result[11] ) );
   NOR2X1 i_31 ( .Y (n_509),
	.B (\ab_result[14] ),
	.A (\ab_result[13] ) );
   NAND3X1 i_110 ( .Y (n_511),
	.C (n_507),
	.B (n_509),
	.A (n_508) );
   NOR2X1 i_32 ( .Y (n_512),
	.B (\ab_result[16] ),
	.A (\ab_result[15] ) );
   NOR2X1 i_33 ( .Y (n_513),
	.B (\ab_result[18] ),
	.A (\ab_result[17] ) );
   NOR4BX1 i_146 ( .Y (n_515),
	.D (n_511),
	.C (\ab_result[16] ),
	.B (\ab_result[15] ),
	.AN (n_513) );
   NOR2X1 i_34 ( .Y (n_516),
	.B (\ab_result[20] ),
	.A (\ab_result[19] ) );
   NOR2X1 i_35 ( .Y (n_517),
	.B (\ab_result[22] ),
	.A (\ab_result[21] ) );
   NAND3X1 i_150 ( .Y (n_519),
	.C (n_515),
	.B (n_517),
	.A (n_516) );
   NOR2X1 i_21 ( .Y (n_520),
	.B (\ab_result[25] ),
	.A (\ab_result[24] ) );
   OR4X1 i_582170 ( .Y (n_522),
	.D (\ab_result[26] ),
	.C (\ab_result[23] ),
	.B (\ab_result[25] ),
	.A (\ab_result[24] ) );
   OR4X1 i_248 ( .Y (n_525),
	.D (\ab_result[30] ),
	.C (\ab_result[29] ),
	.B (\ab_result[28] ),
	.A (\ab_result[27] ) );
   OAI32X1 i_11 ( .Y (n_527),
	.B1 (n_333),
	.B0 (n_334),
	.A2 (n_525),
	.A1 (n_522),
	.A0 (n_519) );
   NOR2X1 i_254 ( .Y (n_528),
	.B (\ab_result[5] ),
	.A (\ab_result[2] ) );
   NAND3X1 i_692179 ( .Y (n_530),
	.C (n_498),
	.B (n_528),
	.A (n_500) );
   NOR4BX1 i_105 ( .Y (n_533),
	.D (n_530),
	.C (\ab_result[9] ),
	.B (\ab_result[6] ),
	.AN (n_504) );
   NOR2X1 i_258 ( .Y (n_534),
	.B (\ab_result[13] ),
	.A (\ab_result[10] ) );
   NAND3X1 i_109 ( .Y (n_536),
	.C (n_533),
	.B (n_534),
	.A (n_508) );
   NOR4BX1 i_145 ( .Y (n_539),
	.D (n_536),
	.C (\ab_result[17] ),
	.B (\ab_result[14] ),
	.AN (n_512) );
   NOR4X1 i_263 ( .Y (n_541),
	.D (\ab_result[21] ),
	.C (\ab_result[18] ),
	.B (\ab_result[20] ),
	.A (\ab_result[19] ) );
   NAND2X1 i_149 ( .Y (n_542),
	.B (n_541),
	.A (n_539) );
   OR4X1 i_572169 ( .Y (n_544),
	.D (\ab_result[25] ),
	.C (\ab_result[24] ),
	.B (\ab_result[23] ),
	.A (\ab_result[22] ) );
   NOR2X1 i_20 ( .Y (n_545),
	.B (\ab_result[27] ),
	.A (\ab_result[26] ) );
   NOR4BX1 i_267 ( .Y (n_548),
	.D (n_544),
	.C (\ab_result[29] ),
	.B (\ab_result[28] ),
	.AN (n_545) );
   AOI31X1 i_12 ( .Y (n_549),
	.B0 (n_268),
	.A2 (n_541),
	.A1 (n_548),
	.A0 (n_539) );
   NAND4X1 i_104 ( .Y (n_552),
	.D (n_504),
	.C (n_501),
	.B (n_500),
	.A (n_499) );
   NOR4BX1 i_108 ( .Y (n_554),
	.D (n_552),
	.C (\ab_result[10] ),
	.B (\ab_result[9] ),
	.AN (n_508) );
   NAND3X1 i_144 ( .Y (n_556),
	.C (n_554),
	.B (n_512),
	.A (n_509) );
   NOR4BX1 i_148 ( .Y (n_558),
	.D (n_556),
	.C (\ab_result[18] ),
	.B (\ab_result[17] ),
	.AN (n_516) );
   NOR4X1 i_562168 ( .Y (n_560),
	.D (\ab_result[24] ),
	.C (\ab_result[23] ),
	.B (\ab_result[22] ),
	.A (\ab_result[21] ) );
   NOR4X1 i_280 ( .Y (n_562),
	.D (\ab_result[28] ),
	.C (\ab_result[25] ),
	.B (\ab_result[27] ),
	.A (\ab_result[26] ) );
   AOI31X1 i_13 ( .Y (n_564),
	.B0 (n_268),
	.A2 (n_562),
	.A1 (n_560),
	.A0 (n_558) );
   NOR3X1 i_287 ( .Y (n_566),
	.C (\ab_result[3] ),
	.B (\ab_result[7] ),
	.A (\ab_result[4] ) );
   NAND3X1 i_712181 ( .Y (n_568),
	.C (n_499),
	.B (n_566),
	.A (n_501) );
   NOR4BX1 i_107 ( .Y (n_571),
	.D (n_568),
	.C (\ab_result[11] ),
	.B (\ab_result[8] ),
	.AN (n_505) );
   NOR2X1 i_291 ( .Y (n_572),
	.B (\ab_result[15] ),
	.A (\ab_result[12] ) );
   NAND3X1 i_111 ( .Y (n_574),
	.C (n_571),
	.B (n_572),
	.A (n_509) );
   NOR4BX1 i_147 ( .Y (n_577),
	.D (n_574),
	.C (\ab_result[19] ),
	.B (\ab_result[16] ),
	.AN (n_513) );
   NOR2X1 i_285 ( .Y (n_578),
	.B (\ab_result[23] ),
	.A (\ab_result[20] ) );
   NAND2X1 i_552167 ( .Y (n_579),
	.B (n_578),
	.A (n_517) );
   NAND2BX1 i_14 ( .Y (n_582),
	.B (n_344),
	.AN (n_268) );
   OAI22X1 i_15 ( .Y (n_583),
	.B1 (n_333),
	.B0 (n_334),
	.A1 (n_522),
	.A0 (n_519) );
   OAI22X1 i_16 ( .Y (n_584),
	.B1 (n_333),
	.B0 (n_334),
	.A1 (n_544),
	.A0 (n_542) );
   AOI21X1 i_17 ( .Y (n_585),
	.B0 (n_268),
	.A1 (n_560),
	.A0 (n_558) );
   AOI31X1 i_18 ( .Y (n_586),
	.B0 (n_268),
	.A2 (n_577),
	.A1 (n_578),
	.A0 (n_517) );
   OAI21XL i_65 ( .Y (n_587),
	.B0 (n_519),
	.A1 (n_333),
	.A0 (n_334) );
   OAI21XL i_66 ( .Y (n_588),
	.B0 (n_542),
	.A1 (n_333),
	.A0 (n_334) );
   NOR2BX1 i_71 ( .Y (n_593),
	.B (n_268),
	.AN (n_556) );
   NOR2BX1 i_72 ( .Y (n_594),
	.B (n_268),
	.AN (n_574) );
   NOR2BX1 i_73 ( .Y (n_595),
	.B (n_268),
	.AN (n_511) );
   NOR2BX1 i_74 ( .Y (n_596),
	.B (n_268),
	.AN (n_536) );
   OAI21XL i_79 ( .Y (n_601),
	.B0 (n_552),
	.A1 (n_333),
	.A0 (n_334) );
   NOR2BX1 i_80 ( .Y (n_602),
	.B (n_268),
	.AN (n_568) );
   NOR2BX1 i_81 ( .Y (n_603),
	.B (n_268),
	.AN (n_503) );
   NOR2BX1 i_82 ( .Y (n_604),
	.B (n_268),
	.AN (n_530) );
   AOI21X1 i_83 ( .Y (n_605),
	.B0 (n_268),
	.A1 (n_500),
	.A0 (n_499) );
   OAI21XL i_86 ( .Y (n_609),
	.B0 (result[0]),
	.A1 (n_333),
	.A0 (n_334) );
   AND4X1 i_248350 ( .Y (\ab_a[15] ),
	.D (n_415),
	.C (op_a[15]),
	.B (n_417),
	.A (n_416) );
   AND4X1 i_248398 ( .Y (\ab_b[15] ),
	.D (n_461),
	.C (op_b[15]),
	.B (n_463),
	.A (n_462) );
   INVX1 i_3316 ( .Y (n_3099),
	.A (n_585) );
   INVX1 i_3317 ( .Y (n_3100),
	.A (n_453) );
   INVX1 i_3318 ( .Y (n_3101),
	.A (n_407) );
   m16x16 M16X16_INST ( .a ({ \ab_a[15] ,
		\ab_a[14] ,
		\ab_a[13] ,
		\ab_a[12] ,
		\ab_a[11] ,
		\ab_a[10] ,
		\ab_a[9] ,
		\ab_a[8] ,
		\ab_a[7] ,
		\ab_a[6] ,
		\ab_a[5] ,
		\ab_a[4] ,
		\ab_a[3] ,
		\ab_a[2] ,
		\ab_a[1] ,
		op_a[0] }),
	.b ({ \ab_b[15] ,
		\ab_b[14] ,
		\ab_b[13] ,
		\ab_b[12] ,
		\ab_b[11] ,
		\ab_b[10] ,
		\ab_b[9] ,
		\ab_b[8] ,
		\ab_b[7] ,
		\ab_b[6] ,
		\ab_b[5] ,
		\ab_b[4] ,
		\ab_b[3] ,
		\ab_b[2] ,
		\ab_b[1] ,
		op_b[0] }),
	.y ({ \ab_result[31] ,
		\ab_result[30] ,
		\ab_result[29] ,
		\ab_result[28] ,
		\ab_result[27] ,
		\ab_result[26] ,
		\ab_result[25] ,
		\ab_result[24] ,
		\ab_result[23] ,
		\ab_result[22] ,
		\ab_result[21] ,
		\ab_result[20] ,
		\ab_result[19] ,
		\ab_result[18] ,
		\ab_result[17] ,
		\ab_result[16] ,
		\ab_result[15] ,
		\ab_result[14] ,
		\ab_result[13] ,
		\ab_result[12] ,
		\ab_result[11] ,
		\ab_result[10] ,
		\ab_result[9] ,
		\ab_result[8] ,
		\ab_result[7] ,
		\ab_result[6] ,
		\ab_result[5] ,
		\ab_result[4] ,
		\ab_result[3] ,
		\ab_result[2] ,
		\ab_result[1] ,
		result[0] }) );
endmodule

module port_bus_mach (
	clk,
	reset,
	read,
	write,
	write_h,
	address,
	data_in,
	data_out,
	pad_data_in,
	pad_data_out,
	addrs_in,
	read_cycle,
	sync,
	go,
	as,
	done,
	scan_en,
	BG_scan_in,
	BG_scan_out );
   input clk;
   input reset;
   output read;
   output write;
   output write_h;
   output [2:0] address;
   input [15:0] data_in;
   output [15:0] data_out;
   input [15:0] pad_data_in;
   output [15:0] pad_data_out;
   input [2:0] addrs_in;
   input read_cycle;
   input sync;
   input go;
   output as;
   output done;
   input scan_en;
   input BG_scan_in;
   output BG_scan_out;

   // Internal wires
   wire [2:0] present_state;
   wire n_6620;
   wire n_6616;
   wire n_6612;
   wire n_6608;
   wire n_6604;
   wire n_6600;
   wire n_6455;
   wire n_6433;
   wire n_6429;
   wire n_6425;
   wire n_6421;
   wire n_6417;
   wire n_6413;
   wire n_6409;
   wire n_6405;
   wire n_6393;
   wire n_11;
   wire n_3051;
   wire n_13;
   wire n_14;
   wire n_15;
   wire \nbus_616[0] ;
   wire n_3052;
   wire FE_OFN136_scan_enI;
   wire n_18;
   wire n_5134;
   wire n_5128;
   wire n_2949;
   wire n_5006;
   wire n_2955;
   wire n_2961;
   wire n_2967;
   wire FE_OFN140_scan_enI;
   wire n_2973;
   wire n_26;
   wire n_21;
   wire n_2979;
   wire FE_OFN141_scan_enI;
   wire n_2985;
   wire n_2991;
   wire FE_OFN12_scan_enI;
   wire n_2997;
   wire n_3003;
   wire n_3009;
   wire n_3015;
   wire n_3021;
   wire n_3027;
   wire n_5042;
   wire FE_OFN15_scan_enI;
   wire n_3033;
   wire n_3039;

   INVX2 i_9768 ( .Y (pad_data_out[2]),
	.A (n_6620) );
   INVXL i_9767 ( .Y (n_6620),
	.A (data_in[2]) );
   INVX2 i_9765 ( .Y (pad_data_out[3]),
	.A (n_6616) );
   INVXL i_9764 ( .Y (n_6616),
	.A (data_in[3]) );
   INVX2 i_9762 ( .Y (pad_data_out[4]),
	.A (n_6612) );
   INVXL i_9761 ( .Y (n_6612),
	.A (data_in[4]) );
   INVX2 i_9759 ( .Y (pad_data_out[5]),
	.A (n_6608) );
   INVXL i_9758 ( .Y (n_6608),
	.A (data_in[5]) );
   INVX2 i_9756 ( .Y (pad_data_out[6]),
	.A (n_6604) );
   INVXL i_9755 ( .Y (n_6604),
	.A (data_in[6]) );
   INVX2 i_9753 ( .Y (pad_data_out[7]),
	.A (n_6600) );
   INVXL i_9752 ( .Y (n_6600),
	.A (data_in[7]) );
   INVX2 i_9644 ( .Y (pad_data_out[1]),
	.A (n_6455) );
   INVXL i_9643 ( .Y (n_6455),
	.A (data_in[1]) );
   INVX2 i_9623 ( .Y (pad_data_out[8]),
	.A (n_6433) );
   INVXL i_9622 ( .Y (n_6433),
	.A (data_in[8]) );
   INVX2 i_9620 ( .Y (pad_data_out[9]),
	.A (n_6429) );
   INVXL i_9619 ( .Y (n_6429),
	.A (data_in[9]) );
   INVX2 i_9617 ( .Y (pad_data_out[10]),
	.A (n_6425) );
   INVXL i_9616 ( .Y (n_6425),
	.A (data_in[10]) );
   INVX2 i_9614 ( .Y (pad_data_out[11]),
	.A (n_6421) );
   INVXL i_9613 ( .Y (n_6421),
	.A (data_in[11]) );
   INVX2 i_9611 ( .Y (pad_data_out[12]),
	.A (n_6417) );
   INVXL i_9610 ( .Y (n_6417),
	.A (data_in[12]) );
   INVX2 i_9608 ( .Y (pad_data_out[13]),
	.A (n_6413) );
   INVXL i_9607 ( .Y (n_6413),
	.A (data_in[13]) );
   INVX2 i_9605 ( .Y (pad_data_out[14]),
	.A (n_6409) );
   INVXL i_9604 ( .Y (n_6409),
	.A (data_in[14]) );
   INVX2 i_9602 ( .Y (pad_data_out[15]),
	.A (n_6405) );
   INVXL i_9601 ( .Y (n_6405),
	.A (data_in[15]) );
   CLKBUFXL i_9600 ( .Y (address[0]),
	.A (addrs_in[0]) );
   CLKBUFXL i_9597 ( .Y (address[1]),
	.A (addrs_in[1]) );
   INVXL i_9593 ( .Y (address[2]),
	.A (n_6393) );
   INVXL i_9592 ( .Y (n_6393),
	.A (addrs_in[2]) );
   CLKBUFX4 i_9504 ( .Y (pad_data_out[0]),
	.A (data_in[0]) );
   AOI211X1 i_11 ( .Y (n_11),
	.C0 (present_state[2]),
	.B0 (present_state[1]),
	.A1 (read_cycle),
	.A0 (go) );
   AOI21X1 i_9 ( .Y (n_13),
	.B0 (n_3051),
	.A1 (present_state[1]),
	.A0 (present_state[0]) );
   NOR4BX1 i_15 ( .Y (n_14),
	.D (present_state[1]),
	.C (present_state[0]),
	.B (read_cycle),
	.AN (go) );
   OR2X1 i_3 ( .Y (n_15),
	.B (n_14),
	.A (n_13) );
   SDFFRHQX1 present_state_reg_0 ( .SI (BG_scan_in),
	.SE (scan_en),
	.RN (n_3052),
	.Q (present_state[0]),
	.D (\nbus_616[0] ),
	.CK (clk) );
   SDFFRHQX1 present_state_reg_1 ( .SI (present_state[0]),
	.SE (FE_OFN136_scan_enI),
	.RN (n_3052),
	.Q (present_state[1]),
	.D (n_18),
	.CK (clk) );
   SDFFRHQX1 present_state_reg_2 ( .SI (present_state[1]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (present_state[2]),
	.D (n_15),
	.CK (clk) );
   SDFFRHQX1 write_reg ( .SI (present_state[2]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (write),
	.D (n_5134),
	.CK (clk) );
   SDFFRHQX1 done_reg ( .SI (write),
	.SE (FE_OFN136_scan_enI),
	.RN (n_3052),
	.Q (done),
	.D (n_5128),
	.CK (clk) );
   SDFFRHQX1 data_out_reg_0 ( .SI (done),
	.SE (scan_en),
	.RN (n_3052),
	.Q (data_out[0]),
	.D (n_2949),
	.CK (clk) );
   MX2X1 i_897 ( .Y (n_2949),
	.S0 (n_5006),
	.B (pad_data_in[0]),
	.A (data_out[0]) );
   SDFFRHQX1 data_out_reg_1 ( .SI (data_out[0]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (data_out[1]),
	.D (n_2955),
	.CK (clk) );
   MX2X1 i_904 ( .Y (n_2955),
	.S0 (n_5006),
	.B (pad_data_in[1]),
	.A (data_out[1]) );
   XOR2X1 i_5 ( .Y (n_18),
	.B (present_state[0]),
	.A (present_state[1]) );
   SDFFRHQX1 data_out_reg_2 ( .SI (data_out[1]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (data_out[2]),
	.D (n_2961),
	.CK (clk) );
   MX2X1 i_911 ( .Y (n_2961),
	.S0 (n_5006),
	.B (pad_data_in[2]),
	.A (data_out[2]) );
   SDFFRHQX1 data_out_reg_3 ( .SI (data_out[2]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (data_out[3]),
	.D (n_2967),
	.CK (clk) );
   MX2X1 i_918 ( .Y (n_2967),
	.S0 (n_5006),
	.B (pad_data_in[3]),
	.A (data_out[3]) );
   SDFFRHQX1 data_out_reg_4 ( .SI (data_out[3]),
	.SE (FE_OFN140_scan_enI),
	.RN (n_3052),
	.Q (data_out[4]),
	.D (n_2973),
	.CK (clk) );
   MX2X1 i_925 ( .Y (n_2973),
	.S0 (n_5006),
	.B (pad_data_in[4]),
	.A (data_out[4]) );
   OR2X1 i_8 ( .Y (n_21),
	.B (n_26),
	.A (n_18) );
   SDFFRHQX1 data_out_reg_5 ( .SI (data_out[4]),
	.SE (FE_OFN140_scan_enI),
	.RN (n_3052),
	.Q (data_out[5]),
	.D (n_2979),
	.CK (clk) );
   MX2X1 i_932 ( .Y (n_2979),
	.S0 (n_5006),
	.B (pad_data_in[5]),
	.A (data_out[5]) );
   SDFFRHQX1 data_out_reg_6 ( .SI (data_out[5]),
	.SE (FE_OFN141_scan_enI),
	.RN (n_3052),
	.Q (data_out[6]),
	.D (n_2985),
	.CK (clk) );
   MX2X1 i_939 ( .Y (n_2985),
	.S0 (n_5006),
	.B (pad_data_in[6]),
	.A (data_out[6]) );
   SDFFRHQX1 data_out_reg_7 ( .SI (data_out[6]),
	.SE (FE_OFN141_scan_enI),
	.RN (n_3052),
	.Q (data_out[7]),
	.D (n_2991),
	.CK (clk) );
   MX2X1 i_946 ( .Y (n_2991),
	.S0 (n_5006),
	.B (pad_data_in[7]),
	.A (data_out[7]) );
   SDFFRHQX1 data_out_reg_8 ( .SI (data_out[7]),
	.SE (FE_OFN12_scan_enI),
	.RN (n_3052),
	.Q (data_out[8]),
	.D (n_2997),
	.CK (clk) );
   MX2X1 i_953 ( .Y (n_2997),
	.S0 (n_5006),
	.B (pad_data_in[8]),
	.A (data_out[8]) );
   SDFFRHQX1 data_out_reg_9 ( .SI (data_out[8]),
	.SE (FE_OFN12_scan_enI),
	.RN (n_3052),
	.Q (data_out[9]),
	.D (n_3003),
	.CK (clk) );
   MX2X1 i_960 ( .Y (n_3003),
	.S0 (n_5006),
	.B (pad_data_in[9]),
	.A (data_out[9]) );
   AOI2BB1X1 i_25 ( .Y (n_26),
	.B0 (present_state[1]),
	.A1N (present_state[2]),
	.A0N (go) );
   SDFFRHQX1 data_out_reg_10 ( .SI (data_out[9]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (data_out[10]),
	.D (n_3009),
	.CK (clk) );
   MX2X1 i_967 ( .Y (n_3009),
	.S0 (n_5006),
	.B (pad_data_in[10]),
	.A (data_out[10]) );
   SDFFRHQX1 data_out_reg_11 ( .SI (data_out[10]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (data_out[11]),
	.D (n_3015),
	.CK (clk) );
   MX2X1 i_974 ( .Y (n_3015),
	.S0 (n_5006),
	.B (pad_data_in[11]),
	.A (data_out[11]) );
   NOR2X1 i_0 ( .Y (n_5134),
	.B (n_3051),
	.A (present_state[1]) );
   SDFFRHQX1 data_out_reg_12 ( .SI (data_out[11]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (data_out[12]),
	.D (n_3021),
	.CK (clk) );
   MX2X1 i_981 ( .Y (n_3021),
	.S0 (n_5006),
	.B (pad_data_in[12]),
	.A (data_out[12]) );
   AND2X1 i_19001 ( .Y (n_5128),
	.B (present_state[0]),
	.A (present_state[1]) );
   SDFFRHQX1 data_out_reg_13 ( .SI (data_out[12]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (data_out[13]),
	.D (n_3027),
	.CK (clk) );
   MX2X1 i_988 ( .Y (n_3027),
	.S0 (n_5006),
	.B (pad_data_in[13]),
	.A (data_out[13]) );
   NOR3BX1 i_2 ( .Y (n_5042),
	.C (present_state[2]),
	.B (present_state[1]),
	.AN (present_state[0]) );
   SDFFRHQX1 data_out_reg_14 ( .SI (data_out[13]),
	.SE (FE_OFN15_scan_enI),
	.RN (n_3052),
	.Q (data_out[14]),
	.D (n_3033),
	.CK (clk) );
   MX2X1 i_995 ( .Y (n_3033),
	.S0 (n_5006),
	.B (pad_data_in[14]),
	.A (data_out[14]) );
   NOR2X1 i_7 ( .Y (\nbus_616[0] ),
	.B (present_state[0]),
	.A (n_11) );
   SDFFRHQX1 data_out_reg_15 ( .SI (data_out[14]),
	.SE (FE_OFN15_scan_enI),
	.RN (n_3052),
	.Q (data_out[15]),
	.D (n_3039),
	.CK (clk) );
   MX2X1 i_1002 ( .Y (n_3039),
	.S0 (n_5006),
	.B (pad_data_in[15]),
	.A (data_out[15]) );
   NOR3BX1 i_10 ( .Y (n_5006),
	.C (present_state[2]),
	.B (present_state[0]),
	.AN (present_state[1]) );
   SDFFRHQX1 read_reg ( .SI (data_out[15]),
	.SE (scan_en),
	.RN (n_3052),
	.Q (read),
	.D (n_5042),
	.CK (clk) );
   SDFFRHQX1 as_reg ( .SI (read),
	.SE (scan_en),
	.RN (n_3052),
	.Q (as),
	.D (n_21),
	.CK (clk) );
   SDFFRHQX1 write_h_reg ( .SI (as),
	.SE (scan_en),
	.RN (n_3052),
	.Q (BG_scan_out),
	.D (n_13),
	.CK (clk) );
   INVX1 i_1069 ( .Y (n_3051),
	.A (present_state[2]) );
   INVX1 i_1070 ( .Y (n_3052),
	.A (reset) );
   BUFX1 FE_OFC141_scan_enI ( .Y (FE_OFN141_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC140_scan_enI ( .Y (FE_OFN140_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC136_scan_enI ( .Y (FE_OFN136_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC15_scan_enI ( .Y (FE_OFN15_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC12_scan_enI ( .Y (FE_OFN12_scan_enI),
	.A (scan_en) );
endmodule

module prog_bus_mach (
	clk,
	reset,
	read,
	write,
	write_h,
	address,
	data_in,
	data_out,
	pad_data_in,
	addrs_in,
	read_cycle,
	sync,
	go,
	as,
	done,
	scan_en,
	BG_scan_in,
	BG_scan_out );
   input clk;
   input reset;
   output read;
   output write;
   output write_h;
   output [8:0] address;
   input [15:0] data_in;
   output [15:0] data_out;
   input [15:0] pad_data_in;
   input [8:0] addrs_in;
   input read_cycle;
   input sync;
   input go;
   output as;
   output done;
   input scan_en;
   input BG_scan_in;
   output BG_scan_out;

   // Internal wires
   wire [2:0] present_state;
   wire n_6491;
   wire n_6487;
   wire n_6483;
   wire n_6479;
   wire n_6475;
   wire n_6471;
   wire n_6467;
   wire n_6463;
   wire n_6459;
   wire n_4835;
   wire n_20;
   wire n_18;
   wire n_17;
   wire \nbus_606[0] ;
   wire n_2937;
   wire n_21;
   wire FE_OFN2_scan_enI;
   wire n_4954;
   wire n_2832;
   wire n_4826;
   wire n_2838;
   wire n_2844;
   wire n_2850;
   wire n_23;
   wire n_4868;
   wire n_2936;
   wire n_2856;
   wire n_2862;
   wire FE_OFN133_scan_enI;
   wire n_2868;
   wire n_2874;
   wire n_25;
   wire n_2880;
   wire n_2886;
   wire n_2892;
   wire n_2898;
   wire n_2904;
   wire n_4862;
   wire n_2910;
   wire n_2916;
   wire n_2922;

   INVXL i_9671 ( .Y (address[0]),
	.A (n_6491) );
   INVXL i_9670 ( .Y (n_6491),
	.A (addrs_in[0]) );
   INVXL i_9668 ( .Y (address[1]),
	.A (n_6487) );
   INVXL i_9667 ( .Y (n_6487),
	.A (addrs_in[1]) );
   INVXL i_9665 ( .Y (address[2]),
	.A (n_6483) );
   INVXL i_9664 ( .Y (n_6483),
	.A (addrs_in[2]) );
   INVXL i_9662 ( .Y (address[3]),
	.A (n_6479) );
   INVXL i_9661 ( .Y (n_6479),
	.A (addrs_in[3]) );
   INVXL i_9659 ( .Y (address[4]),
	.A (n_6475) );
   INVXL i_9658 ( .Y (n_6475),
	.A (addrs_in[4]) );
   INVXL i_9656 ( .Y (address[5]),
	.A (n_6471) );
   INVXL i_9655 ( .Y (n_6471),
	.A (addrs_in[5]) );
   INVXL i_9653 ( .Y (address[6]),
	.A (n_6467) );
   INVXL i_9652 ( .Y (n_6467),
	.A (addrs_in[6]) );
   INVXL i_9650 ( .Y (address[7]),
	.A (n_6463) );
   INVXL i_9649 ( .Y (n_6463),
	.A (addrs_in[7]) );
   INVXL i_9647 ( .Y (address[8]),
	.A (n_6459) );
   INVXL i_9646 ( .Y (n_6459),
	.A (addrs_in[8]) );
   OR3XL i_8 ( .Y (n_17),
	.C (n_18),
	.B (n_20),
	.A (n_4835) );
   SDFFRHQX1 present_state_reg_0 ( .SI (BG_scan_in),
	.SE (scan_en),
	.RN (n_2937),
	.Q (present_state[0]),
	.D (\nbus_606[0] ),
	.CK (clk) );
   SDFFRHQX1 present_state_reg_1 ( .SI (present_state[0]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (present_state[1]),
	.D (n_20),
	.CK (clk) );
   SDFFRHQX1 present_state_reg_2 ( .SI (present_state[1]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (present_state[2]),
	.D (n_21),
	.CK (clk) );
   SDFFRHQX1 write_reg ( .SI (present_state[2]),
	.SE (FE_OFN2_scan_enI),
	.RN (n_2937),
	.Q (write),
	.D (n_4954),
	.CK (clk) );
   SDFFRHQX1 data_out_reg_0 ( .SI (write),
	.SE (FE_OFN2_scan_enI),
	.RN (n_2937),
	.Q (data_out[0]),
	.D (n_2832),
	.CK (clk) );
   MX2X1 i_702 ( .Y (n_2832),
	.S0 (n_4826),
	.B (pad_data_in[0]),
	.A (data_out[0]) );
   NOR2BX1 i_12 ( .Y (n_18),
	.B (present_state[1]),
	.AN (go) );
   SDFFRHQX1 data_out_reg_1 ( .SI (data_out[0]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[1]),
	.D (n_2838),
	.CK (clk) );
   MX2X1 i_709 ( .Y (n_2838),
	.S0 (n_4826),
	.B (pad_data_in[1]),
	.A (data_out[1]) );
   SDFFRHQX1 data_out_reg_2 ( .SI (data_out[1]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[2]),
	.D (n_2844),
	.CK (clk) );
   MX2X1 i_716 ( .Y (n_2844),
	.S0 (n_4826),
	.B (pad_data_in[2]),
	.A (data_out[2]) );
   XOR2X1 i_5 ( .Y (n_20),
	.B (present_state[1]),
	.A (present_state[0]) );
   SDFFRHQX1 data_out_reg_3 ( .SI (data_out[2]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[3]),
	.D (n_2850),
	.CK (clk) );
   MX2X1 i_723 ( .Y (n_2850),
	.S0 (n_4826),
	.B (pad_data_in[3]),
	.A (data_out[3]) );
   OAI32X1 i_3 ( .Y (n_21),
	.B1 (n_2936),
	.B0 (n_4868),
	.A2 (n_23),
	.A1 (present_state[0]),
	.A0 (present_state[1]) );
   SDFFRHQX1 data_out_reg_4 ( .SI (data_out[3]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[4]),
	.D (n_2856),
	.CK (clk) );
   MX2X1 i_730 ( .Y (n_2856),
	.S0 (n_4826),
	.B (pad_data_in[4]),
	.A (data_out[4]) );
   SDFFRHQX1 data_out_reg_5 ( .SI (data_out[4]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[5]),
	.D (n_2862),
	.CK (clk) );
   MX2X1 i_737 ( .Y (n_2862),
	.S0 (n_4826),
	.B (pad_data_in[5]),
	.A (data_out[5]) );
   NAND2BX1 i_25 ( .Y (n_23),
	.B (go),
	.AN (read_cycle) );
   SDFFRHQX1 data_out_reg_6 ( .SI (data_out[5]),
	.SE (FE_OFN133_scan_enI),
	.RN (n_2937),
	.Q (data_out[6]),
	.D (n_2868),
	.CK (clk) );
   MX2X1 i_744 ( .Y (n_2868),
	.S0 (n_4826),
	.B (pad_data_in[6]),
	.A (data_out[6]) );
   SDFFRHQX1 data_out_reg_7 ( .SI (data_out[6]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[7]),
	.D (n_2874),
	.CK (clk) );
   MX2X1 i_751 ( .Y (n_2874),
	.S0 (n_4826),
	.B (pad_data_in[7]),
	.A (data_out[7]) );
   AOI21X1 i_21 ( .Y (n_25),
	.B0 (present_state[1]),
	.A1 (read_cycle),
	.A0 (go) );
   SDFFRHQX1 data_out_reg_8 ( .SI (data_out[7]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[8]),
	.D (n_2880),
	.CK (clk) );
   MX2X1 i_758 ( .Y (n_2880),
	.S0 (n_4826),
	.B (pad_data_in[8]),
	.A (data_out[8]) );
   SDFFRHQX1 data_out_reg_9 ( .SI (data_out[8]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[9]),
	.D (n_2886),
	.CK (clk) );
   MX2X1 i_765 ( .Y (n_2886),
	.S0 (n_4826),
	.B (pad_data_in[9]),
	.A (data_out[9]) );
   SDFFRHQX1 data_out_reg_10 ( .SI (data_out[9]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[10]),
	.D (n_2892),
	.CK (clk) );
   MX2X1 i_772 ( .Y (n_2892),
	.S0 (n_4826),
	.B (pad_data_in[10]),
	.A (data_out[10]) );
   NOR3X1 i_0 ( .Y (n_4954),
	.C (n_2936),
	.B (present_state[0]),
	.A (present_state[1]) );
   SDFFRHQX1 data_out_reg_11 ( .SI (data_out[10]),
	.SE (FE_OFN2_scan_enI),
	.RN (n_2937),
	.Q (data_out[11]),
	.D (n_2898),
	.CK (clk) );
   MX2X1 i_779 ( .Y (n_2898),
	.S0 (n_4826),
	.B (pad_data_in[11]),
	.A (data_out[11]) );
   AND2X1 i_19000 ( .Y (n_4868),
	.B (present_state[0]),
	.A (present_state[1]) );
   SDFFRHQX1 data_out_reg_12 ( .SI (data_out[11]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[12]),
	.D (n_2904),
	.CK (clk) );
   MX2X1 i_786 ( .Y (n_2904),
	.S0 (n_4826),
	.B (pad_data_in[12]),
	.A (data_out[12]) );
   NOR3BX1 i_2 ( .Y (n_4862),
	.C (present_state[2]),
	.B (present_state[1]),
	.AN (present_state[0]) );
   SDFFRHQX1 data_out_reg_13 ( .SI (data_out[12]),
	.SE (FE_OFN2_scan_enI),
	.RN (n_2937),
	.Q (data_out[13]),
	.D (n_2910),
	.CK (clk) );
   MX2X1 i_793 ( .Y (n_2910),
	.S0 (n_4826),
	.B (pad_data_in[13]),
	.A (data_out[13]) );
   AOI21X1 i_7 ( .Y (\nbus_606[0] ),
	.B0 (present_state[0]),
	.A1 (n_2936),
	.A0 (n_25) );
   SDFFRHQX1 data_out_reg_14 ( .SI (data_out[13]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[14]),
	.D (n_2916),
	.CK (clk) );
   MX2X1 i_800 ( .Y (n_2916),
	.S0 (n_4826),
	.B (pad_data_in[14]),
	.A (data_out[14]) );
   NOR2X1 i_9 ( .Y (n_4835),
	.B (n_2936),
	.A (present_state[1]) );
   SDFFRHQX1 data_out_reg_15 ( .SI (data_out[14]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (data_out[15]),
	.D (n_2922),
	.CK (clk) );
   MX2X1 i_807 ( .Y (n_2922),
	.S0 (n_4826),
	.B (pad_data_in[15]),
	.A (data_out[15]) );
   NOR3BX1 i_10 ( .Y (n_4826),
	.C (present_state[2]),
	.B (present_state[0]),
	.AN (present_state[1]) );
   SDFFRHQX1 done_reg ( .SI (data_out[15]),
	.SE (scan_en),
	.RN (n_2937),
	.Q (done),
	.D (n_4868),
	.CK (clk) );
   SDFFRHQX1 read_reg ( .SI (done),
	.SE (FE_OFN133_scan_enI),
	.RN (n_2937),
	.Q (read),
	.D (n_4862),
	.CK (clk) );
   SDFFRHQX1 as_reg ( .SI (read),
	.SE (scan_en),
	.RN (n_2937),
	.Q (as),
	.D (n_17),
	.CK (clk) );
   SDFFRHQX1 write_h_reg ( .SI (as),
	.SE (scan_en),
	.RN (n_2937),
	.Q (BG_scan_out),
	.D (n_4835),
	.CK (clk) );
   INVX1 i_877 ( .Y (n_2936),
	.A (present_state[2]) );
   INVX1 i_878 ( .Y (n_2937),
	.A (reset) );
   BUFX1 FE_OFC133_scan_enI ( .Y (FE_OFN133_scan_enI),
	.A (scan_en) );
   BUFX1 FE_OFC2_scan_enI ( .Y (FE_OFN2_scan_enI),
	.A (scan_en) );
endmodule

module tdsp_core_glue (
	addrs_in,
	data_in,
	p_addrs_in,
	p_data_in,
	port_addrs_in,
	port_data_in,
	ar,
	res_adr,
	res_port_adr,
	se_shift_mdr,
	ze_mdr,
	alu_out,
	go_prog,
	read_prog,
	go_data,
	read_data,
	go_port,
	read_port,
	pc_acc,
	arp,
	ar1,
	ar0,
	dp,
	ir,
	pdr,
	opa,
	opb,
	mdr,
	acc,
	pc,
	data_out,
	p_data_out,
	port_data_out,
	top,
	p,
	alu_cmd,
	sel_op_a,
	sel_op_b,
	dec_go_prog,
	enc_go_prog,
	dec_read_prog,
	enc_read_prog,
	dec_go_data,
	enc_go_data,
	dec_read_data,
	enc_read_data,
	dec_go_port,
	enc_go_port,
	dec_read_port,
	enc_read_port,
	dmov_inc );
   output [7:0] addrs_in;
   output [15:0] data_in;
   output [8:0] p_addrs_in;
   output [15:0] p_data_in;
   output [2:0] port_addrs_in;
   output [15:0] port_data_in;
   output [15:0] ar;
   output [7:0] res_adr;
   output [7:0] res_port_adr;
   output [31:0] se_shift_mdr;
   output [31:0] ze_mdr;
   output [15:0] alu_out;
   output go_prog;
   output read_prog;
   output go_data;
   output read_data;
   output go_port;
   output read_port;
   input pc_acc;
   input arp;
   input [15:0] ar1;
   input [15:0] ar0;
   input dp;
   input [15:0] ir;
   output [15:0] pdr;
   output [31:0] opa;
   output [31:0] opb;
   output [15:0] mdr;
   input [32:0] acc;
   input [15:0] pc;
   input [15:0] data_out;
   input [15:0] p_data_out;
   input [15:0] port_data_out;
   input [15:0] top;
   input [31:0] p;
   input [3:0] alu_cmd;
   input [2:0] sel_op_a;
   input [2:0] sel_op_b;
   input dec_go_prog;
   input enc_go_prog;
   input dec_read_prog;
   input enc_read_prog;
   input dec_go_data;
   input enc_go_data;
   input dec_read_data;
   input enc_read_data;
   input dec_go_port;
   input enc_go_port;
   input dec_read_port;
   input enc_read_port;
   input dmov_inc;

   // Internal wires
   wire n_6563;
   wire n_6559;
   wire n_6555;
   wire n_6551;
   wire n_6547;
   wire n_6543;
   wire n_6539;
   wire n_6535;
   wire n_6531;
   wire n_6527;
   wire n_6523;
   wire n_6519;
   wire n_6515;
   wire n_6511;
   wire n_6507;
   wire n_6503;
   wire n_6499;
   wire n_6495;
   wire FE_OFN94_n_1023;
   wire n_1026;
   wire n_1015;
   wire n_1100;
   wire n_1045;
   wire FE_OFN92_n_1037;
   wire n_952;
   wire n_1097;
   wire n_557;
   wire n_1049;
   wire n_571;
   wire n_1086;
   wire n_563;
   wire n_1050;
   wire n_1096;
   wire FE_OFN93_n_1035;
   wire n_1093;
   wire n_1092;
   wire n_962;
   wire n_1089;
   wire n_560;
   wire n_580;
   wire n_566;
   wire n_1088;
   wire n_1084;
   wire n_1083;
   wire n_1079;
   wire n_1080;
   wire n_1069;
   wire n_570;
   wire n_1077;
   wire n_1078;
   wire n_1040;
   wire n_1042;
   wire n_1075;
   wire n_1074;
   wire n_1070;
   wire n_1071;
   wire n_579;
   wire n_1038;
   wire n_1067;
   wire n_1068;
   wire n_1065;
   wire n_1064;
   wire n_1046;
   wire n_4527;
   wire n_1061;
   wire n_997;
   wire n_1059;
   wire n_1056;
   wire n_1055;
   wire n_4526;
   wire n_1052;
   wire n_1048;
   wire n_1013;
   wire n_1021;
   wire n_1008;
   wire n_1044;
   wire n_452;
   wire n_1041;
   wire n_4506;
   wire n_4525;
   wire n_1039;
   wire n_1027;
   wire n_1037;
   wire n_1016;
   wire n_1030;
   wire n_1011;
   wire n_1035;
   wire n_1031;
   wire n_1020;
   wire n_1023;
   wire n_1017;
   wire n_4508;
   wire n_578;
   wire n_569;
   wire n_942;
   wire n_932;
   wire n_922;
   wire n_912;
   wire n_554;
   wire n_902;
   wire n_551;
   wire n_892;
   wire n_863;
   wire n_852;
   wire n_851;
   wire n_850;
   wire n_1215;
   wire n_832;
   wire n_1213;
   wire n_808;
   wire n_1220;
   wire n_807;
   wire n_799;
   wire n_791;
   wire n_783;
   wire n_1221;
   wire n_775;
   wire n_446;
   wire n_4507;
   wire n_758;
   wire n_438;
   wire n_4511;
   wire n_757;
   wire n_4504;
   wire n_719;
   wire n_1314;
   wire n_1218;
   wire n_701;
   wire n_672;
   wire n_667;
   wire n_1308;
   wire n_660;
   wire n_657;
   wire n_1359;
   wire n_604;
   wire n_600;
   wire n_592;
   wire n_548;
   wire n_545;
   wire n_542;
   wire n_539;
   wire n_1208;
   wire n_1194;
   wire n_489;
   wire n_1207;
   wire n_1195;
   wire n_487;
   wire n_1206;
   wire n_1196;
   wire n_485;
   wire n_1205;
   wire n_1197;
   wire n_483;
   wire n_1204;
   wire n_1198;
   wire n_482;
   wire n_1210;
   wire n_1199;
   wire n_480;
   wire n_1209;
   wire n_1201;
   wire n_478;
   wire n_456;
   wire n_449;
   wire n_447;
   wire n_1228;
   wire n_1227;
   wire n_1232;
   wire n_1231;
   wire n_445;
   wire n_1236;
   wire n_1235;
   wire n_444;
   wire n_4510;
   wire n_443;
   wire n_1247;
   wire n_1246;
   wire n_442;
   wire n_1252;
   wire n_1251;
   wire n_441;
   wire n_1257;
   wire n_1256;
   wire n_440;
   wire n_1264;
   wire n_1263;
   wire n_439;
   wire n_1270;
   wire n_1269;
   wire n_1276;
   wire n_1275;
   wire n_437;
   wire n_1282;
   wire n_1281;
   wire n_436;
   wire n_1289;
   wire n_1288;
   wire n_435;
   wire n_432;
   wire n_1294;
   wire n_430;
   wire n_428;
   wire n_4520;
   wire n_410;
   wire n_402;
   wire n_1101;
   wire n_1104;
   wire n_1105;
   wire n_1108;
   wire n_1109;
   wire n_1112;
   wire n_1113;
   wire n_1116;
   wire n_1117;
   wire n_1120;
   wire n_1121;
   wire n_1124;
   wire n_1125;
   wire n_1128;
   wire n_1129;
   wire n_1132;
   wire n_1133;
   wire n_1136;
   wire n_1137;
   wire n_1140;
   wire n_1141;
   wire n_1144;
   wire n_1145;
   wire n_1148;
   wire n_1149;
   wire n_1152;
   wire n_4514;
   wire n_1153;
   wire n_1154;
   wire n_1155;
   wire n_1156;
   wire n_1159;
   wire n_1160;
   wire n_1163;
   wire n_1164;
   wire n_1165;
   wire n_1166;
   wire n_1169;
   wire n_1170;
   wire n_1172;
   wire n_1173;
   wire n_1174;
   wire n_1176;
   wire n_4513;
   wire n_1179;
   wire n_1181;
   wire n_1187;
   wire n_1188;
   wire n_1190;
   wire n_1192;
   wire ar_36576;
   wire n_4524;
   wire ar_26577;
   wire n_4523;
   wire ar_06579;
   wire n_4521;
   wire n_1200;
   wire ar_16578;
   wire n_4522;
   wire n_1211;
   wire n_1214;
   wire n_1216;
   wire n_1217;
   wire n_4496;
   wire n_1219;
   wire n_1222;
   wire n_1223;
   wire n_1226;
   wire n_1229;
   wire n_1230;
   wire n_1233;
   wire n_1234;
   wire n_1237;
   wire n_1239;
   wire n_1241;
   wire n_4509;
   wire n_1243;
   wire n_1244;
   wire n_1249;
   wire n_1254;
   wire n_1258;
   wire n_1260;
   wire n_1261;
   wire n_4498;
   wire n_1266;
   wire n_1267;
   wire n_1272;
   wire n_1273;
   wire n_1278;
   wire n_1279;
   wire n_1283;
   wire n_4499;
   wire n_4497;
   wire n_1285;
   wire n_1287;
   wire n_4500;
   wire n_1291;
   wire n_1293;
   wire n_4505;
   wire n_1295;
   wire n_1296;
   wire n_1298;
   wire n_1299;
   wire n_1300;
   wire n_4502;
   wire n_1303;
   wire n_1304;
   wire n_1306;
   wire n_1309;
   wire n_1310;
   wire n_1312;
   wire n_1315;
   wire n_1316;
   wire n_1318;
   wire n_1320;
   wire n_1323;
   wire n_1324;
   wire n_1327;
   wire n_1328;
   wire n_1331;
   wire n_1332;
   wire n_1335;
   wire n_1336;
   wire n_1338;
   wire n_1339;
   wire n_1341;
   wire n_1342;
   wire n_1343;
   wire n_1344;
   wire n_1345;
   wire n_1347;
   wire n_1349;
   wire n_1351;
   wire n_1352;
   wire n_1353;
   wire n_1355;
   wire n_1357;
   wire n_1358;
   wire n_1360;
   wire n_1361;
   wire n_1362;
   wire n_1363;
   wire n_1364;
   wire n_1365;
   wire n_1366;
   wire n_1367;
   wire n_1368;
   wire n_1369;
   wire n_1370;
   wire n_1371;
   wire n_1372;
   wire n_1373;
   wire n_1374;
   wire n_1375;
   wire n_1376;
   wire n_1378;
   wire n_1380;
   wire n_1381;
   wire n_1382;
   wire n_1384;
   wire opb_316580;
   wire n_4512;
   wire n_4501;
   wire n_4503;

   INVX2 i_9833 ( .Y (mdr[0]),
	.A (n_6563) );
   INVXL i_9829 ( .Y (mdr[1]),
	.A (n_6559) );
   INVXL i_9825 ( .Y (mdr[2]),
	.A (n_6555) );
   INVXL i_9821 ( .Y (mdr[3]),
	.A (n_6551) );
   INVXL i_9817 ( .Y (mdr[4]),
	.A (n_6547) );
   INVXL i_9813 ( .Y (mdr[5]),
	.A (n_6543) );
   INVX2 i_9809 ( .Y (mdr[6]),
	.A (n_6539) );
   INVXL i_9805 ( .Y (mdr[7]),
	.A (n_6535) );
   INVXL i_9801 ( .Y (mdr[8]),
	.A (n_6531) );
   INVXL i_9797 ( .Y (mdr[9]),
	.A (n_6527) );
   INVXL i_9793 ( .Y (mdr[10]),
	.A (n_6523) );
   INVXL i_9789 ( .Y (mdr[11]),
	.A (n_6519) );
   INVXL i_9785 ( .Y (mdr[12]),
	.A (n_6515) );
   INVXL i_9781 ( .Y (mdr[13]),
	.A (n_6511) );
   INVXL i_9777 ( .Y (mdr[14]),
	.A (n_6507) );
   INVXL i_9773 ( .Y (mdr[15]),
	.A (n_6503) );
   INVXL i_9725 ( .Y (port_data_in[0]),
	.A (n_6563) );
   INVXL i_9724 ( .Y (n_6563),
	.A (data_out[0]) );
   INVXL i_9722 ( .Y (port_data_in[1]),
	.A (n_6559) );
   INVXL i_9721 ( .Y (n_6559),
	.A (data_out[1]) );
   INVXL i_9719 ( .Y (port_data_in[2]),
	.A (n_6555) );
   INVXL i_9718 ( .Y (n_6555),
	.A (data_out[2]) );
   INVXL i_9716 ( .Y (port_data_in[3]),
	.A (n_6551) );
   INVXL i_9715 ( .Y (n_6551),
	.A (data_out[3]) );
   INVXL i_9713 ( .Y (port_data_in[4]),
	.A (n_6547) );
   INVXL i_9712 ( .Y (n_6547),
	.A (data_out[4]) );
   INVXL i_9710 ( .Y (port_data_in[5]),
	.A (n_6543) );
   INVXL i_9709 ( .Y (n_6543),
	.A (data_out[5]) );
   INVXL i_9707 ( .Y (port_data_in[6]),
	.A (n_6539) );
   INVXL i_9706 ( .Y (n_6539),
	.A (data_out[6]) );
   INVXL i_9704 ( .Y (port_data_in[7]),
	.A (n_6535) );
   INVXL i_9703 ( .Y (n_6535),
	.A (data_out[7]) );
   INVXL i_9701 ( .Y (port_data_in[8]),
	.A (n_6531) );
   INVXL i_9700 ( .Y (n_6531),
	.A (data_out[8]) );
   INVXL i_9698 ( .Y (port_data_in[9]),
	.A (n_6527) );
   INVXL i_9697 ( .Y (n_6527),
	.A (data_out[9]) );
   INVXL i_9695 ( .Y (port_data_in[10]),
	.A (n_6523) );
   INVXL i_9694 ( .Y (n_6523),
	.A (data_out[10]) );
   INVXL i_9692 ( .Y (port_data_in[11]),
	.A (n_6519) );
   INVXL i_9691 ( .Y (n_6519),
	.A (data_out[11]) );
   INVXL i_9689 ( .Y (port_data_in[12]),
	.A (n_6515) );
   INVXL i_9688 ( .Y (n_6515),
	.A (data_out[12]) );
   INVXL i_9686 ( .Y (port_data_in[13]),
	.A (n_6511) );
   INVXL i_9685 ( .Y (n_6511),
	.A (data_out[13]) );
   INVXL i_9683 ( .Y (port_data_in[14]),
	.A (n_6507) );
   INVXL i_9682 ( .Y (n_6507),
	.A (data_out[14]) );
   INVXL i_9680 ( .Y (port_data_in[15]),
	.A (n_6503) );
   INVXL i_9679 ( .Y (n_6503),
	.A (data_out[15]) );
   INVX1 i_9677 ( .Y (port_addrs_in[0]),
	.A (n_6499) );
   INVXL i_9676 ( .Y (n_6499),
	.A (ir[8]) );
   INVX1 i_9674 ( .Y (port_addrs_in[2]),
	.A (n_6495) );
   INVXL i_9673 ( .Y (n_6495),
	.A (ir[10]) );
   BUFX3 i_9483 ( .Y (port_addrs_in[1]),
	.A (ir[9]) );
   AOI222X1 i_935 ( .Y (n_1100),
	.C1 (n_1015),
	.C0 (port_data_out[5]),
	.B1 (n_1026),
	.B0 (ar1[5]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[5]) );
   AOI31X1 i_937 ( .Y (n_1097),
	.B0 (n_952),
	.A2 (acc[5]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   OAI222XL i_939 ( .Y (n_1096),
	.C1 (n_1050),
	.C0 (n_563),
	.B1 (n_1086),
	.B0 (n_571),
	.A1 (n_1049),
	.A0 (n_557) );
   AOI22X1 i_941 ( .Y (n_1093),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[4]),
	.A1 (dmov_inc),
	.A0 (mdr[4]) );
   AOI222X1 i_943 ( .Y (n_1092),
	.C1 (n_1015),
	.C0 (port_data_out[4]),
	.B1 (n_1026),
	.B0 (ar1[4]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[4]) );
   AOI31X1 i_945 ( .Y (n_1089),
	.B0 (n_962),
	.A2 (acc[4]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   OAI222XL i_947 ( .Y (n_1088),
	.C1 (n_1050),
	.C0 (n_566),
	.B1 (n_1086),
	.B0 (n_580),
	.A1 (n_1049),
	.A0 (n_560) );
   NAND3X1 i_33 ( .Y (n_1086),
	.C (port_addrs_in[1]),
	.B (FE_OFN92_n_1037),
	.A (port_addrs_in[2]) );
   AOI22X1 i_949 ( .Y (n_1084),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[3]),
	.A1 (dmov_inc),
	.A0 (mdr[3]) );
   AOI222X1 i_951 ( .Y (n_1083),
	.C1 (n_1015),
	.C0 (port_data_out[3]),
	.B1 (n_1026),
	.B0 (ar1[3]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[3]) );
   AOI31X1 i_954 ( .Y (n_1080),
	.B0 (n_1079),
	.A2 (acc[3]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   OAI22X1 i_953 ( .Y (n_1079),
	.B1 (n_1050),
	.B0 (n_570),
	.A1 (n_1069),
	.A0 (n_571) );
   OAI21XL i_956 ( .Y (n_1078),
	.B0 (n_1077),
	.A1 (n_1049),
	.A0 (n_563) );
   AOI22X1 i_955 ( .Y (n_1077),
	.B1 (n_1042),
	.B0 (acc[12]),
	.A1 (n_1040),
	.A0 (acc[13]) );
   AOI22X1 i_958 ( .Y (n_1075),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[2]),
	.A1 (dmov_inc),
	.A0 (mdr[2]) );
   AOI222X1 i_960 ( .Y (n_1074),
	.C1 (n_1015),
	.C0 (port_data_out[2]),
	.B1 (n_1026),
	.B0 (ar1[2]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[2]) );
   AOI31X1 i_963 ( .Y (n_1071),
	.B0 (n_1070),
	.A2 (acc[2]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   OAI22X1 i_962 ( .Y (n_1070),
	.B1 (n_1050),
	.B0 (n_579),
	.A1 (n_1069),
	.A0 (n_580) );
   OR2X1 i_30 ( .Y (n_1069),
	.B (n_1038),
	.A (port_addrs_in[1]) );
   OAI21XL i_965 ( .Y (n_1068),
	.B0 (n_1067),
	.A1 (n_1049),
	.A0 (n_566) );
   AOI22X1 i_964 ( .Y (n_1067),
	.B1 (n_1042),
	.B0 (acc[11]),
	.A1 (n_1040),
	.A0 (acc[12]) );
   AOI22X1 i_967 ( .Y (n_1065),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[1]),
	.A1 (dmov_inc),
	.A0 (mdr[1]) );
   AOI222X1 i_969 ( .Y (n_1064),
	.C1 (n_1015),
	.C0 (port_data_out[1]),
	.B1 (n_1026),
	.B0 (ar1[1]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[1]) );
   OAI222XL i_972 ( .Y (n_1061),
	.C1 (n_4527),
	.C0 (n_1046),
	.B1 (n_1049),
	.B0 (n_570),
	.A1 (n_1050),
	.A0 (n_571) );
   AOI221X1 i_974 ( .Y (n_1059),
	.C0 (n_997),
	.B1 (n_1040),
	.B0 (acc[11]),
	.A1 (n_1042),
	.A0 (acc[10]) );
   AOI22X1 i_976 ( .Y (n_1056),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[0]),
	.A1 (mdr[0]),
	.A0 (dmov_inc) );
   AOI222X1 i_978 ( .Y (n_1055),
	.C1 (n_1015),
	.C0 (port_data_out[0]),
	.B1 (n_1026),
	.B0 (ar1[0]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[0]) );
   OAI222XL i_981 ( .Y (n_1052),
	.C1 (n_4526),
	.C0 (n_1046),
	.B1 (n_1049),
	.B0 (n_579),
	.A1 (n_1050),
	.A0 (n_580) );
   NAND2X1 i_31 ( .Y (n_1050),
	.B (n_1048),
	.A (port_addrs_in[1]) );
   NAND2BX1 i_32 ( .Y (n_1049),
	.B (n_1048),
	.AN (port_addrs_in[1]) );
   NOR3BX1 i_4 ( .Y (n_1048),
	.C (n_1045),
	.B (port_addrs_in[2]),
	.AN (FE_OFN92_n_1037) );
   NAND2X1 i_9 ( .Y (n_1046),
	.B (FE_OFN92_n_1037),
	.A (n_1045) );
   NOR2X1 i_60 ( .Y (n_1045),
	.B (n_1021),
	.A (n_1013) );
   AOI221X1 i_983 ( .Y (n_1044),
	.C0 (n_1008),
	.B1 (n_1040),
	.B0 (acc[10]),
	.A1 (n_1042),
	.A0 (acc[9]) );
   NOR2X1 i_65 ( .Y (n_1042),
	.B (n_1038),
	.A (n_452) );
   NOR2X2 i_21 ( .Y (n_1041),
	.B (port_addrs_in[1]),
	.A (ir[8]) );
   NOR2X1 i_62 ( .Y (n_1040),
	.B (n_1038),
	.A (n_4506) );
   NOR2X1 i_20 ( .Y (n_1039),
	.B (n_4525),
	.A (ir[8]) );
   NAND2X1 i_6 ( .Y (n_1038),
	.B (FE_OFN92_n_1037),
	.A (port_addrs_in[2]) );
   NOR4BX1 i_5419 ( .Y (n_1037),
	.D (n_1015),
	.C (FE_OFN93_n_1035),
	.B (dmov_inc),
	.AN (n_1027) );
   NOR4BX1 i_5409 ( .Y (n_1035),
	.D (n_1011),
	.C (n_1030),
	.B (n_1016),
	.AN (port_addrs_in[2]) );
   AND2X1 i_22 ( .Y (n_1031),
	.B (n_4525),
	.A (ir[8]) );
   NAND3BX1 i_992 ( .Y (n_1030),
	.C (ir[14]),
	.B (ir[15]),
	.AN (ir[12]) );
   NOR2X1 i_987 ( .Y (n_1027),
	.B (FE_OFN94_n_1023),
	.A (n_1026) );
   NOR4BBX2 i_5418 ( .Y (n_1026),
	.D (ir[14]),
	.C (n_1016),
	.BN (ir[8]),
	.AN (n_1020) );
   NOR4BX1 i_5415 ( .Y (n_1023),
	.D (n_1016),
	.C (ir[14]),
	.B (ir[8]),
	.AN (n_1020) );
   NAND2BX1 i_58 ( .Y (n_1021),
	.B (n_1020),
	.AN (ir[8]) );
   NOR4BX1 i_16 ( .Y (n_1020),
	.D (n_1017),
	.C (ir[15]),
	.B (port_addrs_in[2]),
	.AN (n_4525) );
   NAND2BX1 i_999 ( .Y (n_1017),
	.B (ir[12]),
	.AN (ir[11]) );
   NAND2BX1 i_70 ( .Y (n_1016),
	.B (ir[13]),
	.AN (dmov_inc) );
   NOR4X2 i_5412 ( .Y (n_1015),
	.D (dmov_inc),
	.C (ir[12]),
	.B (n_1013),
	.A (ir[15]) );
   NAND2BX1 i_57 ( .Y (n_1013),
	.B (ir[14]),
	.AN (ir[13]) );
   MXI2X1 i_53 ( .Y (n_1011),
	.S0 (ir[11]),
	.B (n_1031),
	.A (n_4508) );
   NOR2X1 i_666 ( .Y (n_1008),
	.B (n_1038),
	.A (n_578) );
   NOR2X1 i_649 ( .Y (n_997),
	.B (n_1038),
	.A (n_569) );
   NOR2X1 i_614 ( .Y (n_962),
	.B (n_1069),
	.A (n_579) );
   NOR2X1 i_602 ( .Y (n_952),
	.B (n_1069),
	.A (n_570) );
   NOR2X1 i_590 ( .Y (n_942),
	.B (n_1069),
	.A (n_566) );
   NOR2X1 i_569 ( .Y (n_932),
	.B (n_1069),
	.A (n_563) );
   NOR2X1 i_557 ( .Y (n_922),
	.B (n_1069),
	.A (n_560) );
   NOR2X1 i_513 ( .Y (n_912),
	.B (n_1069),
	.A (n_557) );
   NOR2X1 i_501 ( .Y (n_902),
	.B (n_1069),
	.A (n_554) );
   NOR2X1 i_489 ( .Y (n_892),
	.B (n_1069),
	.A (n_551) );
   NAND3XL i_453 ( .Y (n_863),
	.C (acc[30]),
	.B (n_1048),
	.A (n_1041) );
   NAND3X1 i_442 ( .Y (n_852),
	.C (acc[30]),
	.B (n_1048),
	.A (n_1031) );
   NAND3X1 i_441 ( .Y (n_851),
	.C (acc[31]),
	.B (n_1048),
	.A (n_1041) );
   NAND3BX1 i_440 ( .Y (n_850),
	.C (n_1048),
	.B (acc[29]),
	.AN (n_4506) );
   NOR2BX1 i_581 ( .Y (p_addrs_in[8]),
	.B (pc_acc),
	.AN (pc[8]) );
   NAND2X1 i_343 ( .Y (n_832),
	.B (n_1215),
	.A (mdr[12]) );
   NAND2X1 i_323 ( .Y (n_808),
	.B (n_1213),
	.A (p[25]) );
   NAND2X1 i_13 ( .Y (n_807),
	.B (n_1220),
	.A (mdr[15]) );
   NAND2X1 i_315 ( .Y (n_799),
	.B (n_1213),
	.A (p[24]) );
   NAND2X1 i_307 ( .Y (n_791),
	.B (n_1213),
	.A (p[23]) );
   NAND2X1 i_299 ( .Y (n_783),
	.B (n_1213),
	.A (p[22]) );
   NAND2BX1 i_66 ( .Y (n_775),
	.B (n_1220),
	.AN (n_1221) );
   AND2X1 i_270 ( .Y (n_758),
	.B (n_4507),
	.A (n_446) );
   AND2X1 i_269 ( .Y (n_757),
	.B (n_4511),
	.A (n_438) );
   NAND2X1 i_63 ( .Y (n_719),
	.B (n_4504),
	.A (ir[12]) );
   NOR2X1 i_208 ( .Y (n_701),
	.B (n_1218),
	.A (n_1314) );
   NAND2X1 i_181 ( .Y (n_672),
	.B (n_4504),
	.A (ir[7]) );
   NAND2X1 i_176 ( .Y (n_667),
	.B (n_4504),
	.A (ir[6]) );
   NAND2X1 i_169 ( .Y (n_660),
	.B (n_4507),
	.A (n_1308) );
   NAND2X1 i_166 ( .Y (n_657),
	.B (n_4504),
	.A (ir[4]) );
   NAND2X1 i_89 ( .Y (n_604),
	.B (n_1359),
	.A (top[3]) );
   NAND2X1 i_85 ( .Y (n_600),
	.B (n_1359),
	.A (top[2]) );
   NAND2X1 i_77 ( .Y (n_592),
	.B (n_1359),
	.A (top[0]) );
   MXI2X1 i_152250 ( .Y (n_580),
	.S0 (port_addrs_in[0]),
	.B (acc[13]),
	.A (acc[14]) );
   MXI2X1 i_172252 ( .Y (n_579),
	.S0 (port_addrs_in[0]),
	.B (acc[15]),
	.A (acc[16]) );
   AOI22X1 i_72 ( .Y (n_578),
	.B1 (n_1031),
	.B0 (acc[11]),
	.A1 (n_1041),
	.A0 (acc[12]) );
   MXI2X1 i_162251 ( .Y (n_571),
	.S0 (port_addrs_in[0]),
	.B (acc[14]),
	.A (acc[15]) );
   MXI2X1 i_182253 ( .Y (n_570),
	.S0 (port_addrs_in[0]),
	.B (acc[16]),
	.A (acc[17]) );
   AOI22X1 i_73 ( .Y (n_569),
	.B1 (n_1031),
	.B0 (acc[12]),
	.A1 (n_1041),
	.A0 (acc[13]) );
   MXI2X1 i_192254 ( .Y (n_566),
	.S0 (port_addrs_in[0]),
	.B (acc[17]),
	.A (acc[18]) );
   MXI2X1 i_202255 ( .Y (n_563),
	.S0 (port_addrs_in[0]),
	.B (acc[18]),
	.A (acc[19]) );
   MXI2X1 i_212256 ( .Y (n_560),
	.S0 (port_addrs_in[0]),
	.B (acc[19]),
	.A (acc[20]) );
   MXI2X1 i_222257 ( .Y (n_557),
	.S0 (port_addrs_in[0]),
	.B (acc[20]),
	.A (acc[21]) );
   MXI2X1 i_23 ( .Y (n_554),
	.S0 (port_addrs_in[0]),
	.B (acc[21]),
	.A (acc[22]) );
   MXI2X1 i_242258 ( .Y (n_551),
	.S0 (port_addrs_in[0]),
	.B (acc[22]),
	.A (acc[23]) );
   MXI2X1 i_252259 ( .Y (n_548),
	.S0 (ir[8]),
	.B (acc[23]),
	.A (acc[24]) );
   MXI2X1 i_262260 ( .Y (n_545),
	.S0 (ir[8]),
	.B (acc[24]),
	.A (acc[25]) );
   MXI2X1 i_272261 ( .Y (n_542),
	.S0 (port_addrs_in[0]),
	.B (acc[25]),
	.A (acc[26]) );
   MXI2X1 i_282262 ( .Y (n_539),
	.S0 (port_addrs_in[0]),
	.B (acc[26]),
	.A (acc[27]) );
   NAND2X1 i_390 ( .Y (n_489),
	.B (n_1194),
	.A (n_1208) );
   NAND2X1 i_388 ( .Y (n_487),
	.B (n_1195),
	.A (n_1207) );
   NAND2X1 i_386 ( .Y (n_485),
	.B (n_1196),
	.A (n_1206) );
   NAND2X1 i_384 ( .Y (n_483),
	.B (n_1197),
	.A (n_1205) );
   NAND2X1 i_383 ( .Y (n_482),
	.B (n_1198),
	.A (n_1204) );
   NAND2X1 i_381 ( .Y (n_480),
	.B (n_1199),
	.A (n_1210) );
   NAND2X1 i_379 ( .Y (n_478),
	.B (n_1201),
	.A (n_1209) );
   AOI21X1 i_74 ( .Y (n_456),
	.B0 (sel_op_b[2]),
	.A1 (sel_op_b[1]),
	.A0 (sel_op_b[0]) );
   NAND2X1 i_75 ( .Y (n_452),
	.B (port_addrs_in[1]),
	.A (ir[8]) );
   AOI22X1 i_51 ( .Y (n_449),
	.B1 (n_452),
	.B0 (mdr[15]),
	.A1 (n_4508),
	.A0 (mdr[14]) );
   AOI222X1 i_50 ( .Y (n_447),
	.C1 (n_4525),
	.C0 (mdr[15]),
	.B1 (n_1039),
	.B0 (mdr[14]),
	.A1 (n_4508),
	.A0 (mdr[13]) );
   NAND2X1 i_49 ( .Y (n_446),
	.B (n_1227),
	.A (n_1228) );
   NAND2X1 i_48 ( .Y (n_445),
	.B (n_1231),
	.A (n_1232) );
   NAND2X1 i_47 ( .Y (n_444),
	.B (n_1235),
	.A (n_1236) );
   AOI221XL i_46 ( .Y (n_443),
	.C0 (n_4510),
	.B1 (n_1039),
	.B0 (mdr[10]),
	.A1 (n_4508),
	.A0 (mdr[9]) );
   NAND2X1 i_45 ( .Y (n_442),
	.B (n_1246),
	.A (n_1247) );
   NAND2X1 i_44 ( .Y (n_441),
	.B (n_1251),
	.A (n_1252) );
   NAND2X1 i_43 ( .Y (n_440),
	.B (n_1256),
	.A (n_1257) );
   NAND2X1 i_42 ( .Y (n_439),
	.B (n_1263),
	.A (n_1264) );
   NAND2X1 i_41 ( .Y (n_438),
	.B (n_1269),
	.A (n_1270) );
   NAND2X1 i_40 ( .Y (n_437),
	.B (n_1275),
	.A (n_1276) );
   NAND2X1 i_39 ( .Y (n_436),
	.B (n_1281),
	.A (n_1282) );
   NAND2X1 i_38 ( .Y (n_435),
	.B (n_1288),
	.A (n_1289) );
   MXI2X1 i_22222 ( .Y (n_432),
	.S0 (port_addrs_in[0]),
	.B (mdr[0]),
	.A (mdr[1]) );
   OAI21XL i_37 ( .Y (n_430),
	.B0 (n_1294),
	.A1 (n_4525),
	.A0 (n_432) );
   AOI222X1 i_36 ( .Y (n_428),
	.C1 (n_1039),
	.C0 (mdr[0]),
	.B1 (n_1031),
	.B0 (mdr[1]),
	.A1 (n_1041),
	.A0 (mdr[2]) );
   OAI21XL i_09007 ( .Y (n_410),
	.B0 (sel_op_a[0]),
	.A1 (n_4520),
	.A0 (sel_op_a[1]) );
   NAND2X1 i_7 ( .Y (n_402),
	.B (n_410),
	.A (mdr[15]) );
   AOI22X1 i_933 ( .Y (n_1101),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[5]),
	.A1 (dmov_inc),
	.A0 (mdr[5]) );
   OAI222XL i_931 ( .Y (n_1104),
	.C1 (n_1050),
	.C0 (n_560),
	.B1 (n_1086),
	.B0 (n_579),
	.A1 (n_1049),
	.A0 (n_554) );
   AOI31X1 i_929 ( .Y (n_1105),
	.B0 (n_942),
	.A2 (acc[6]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   AOI222X1 i_927 ( .Y (n_1108),
	.C1 (n_1015),
	.C0 (port_data_out[6]),
	.B1 (n_1026),
	.B0 (ar1[6]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[6]) );
   AOI22X1 i_925 ( .Y (n_1109),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[6]),
	.A1 (dmov_inc),
	.A0 (mdr[6]) );
   OAI222XL i_923 ( .Y (n_1112),
	.C1 (n_1050),
	.C0 (n_557),
	.B1 (n_1086),
	.B0 (n_570),
	.A1 (n_1049),
	.A0 (n_551) );
   AOI31X1 i_921 ( .Y (n_1113),
	.B0 (n_932),
	.A2 (acc[7]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   AOI222X1 i_919 ( .Y (n_1116),
	.C1 (n_1015),
	.C0 (port_data_out[7]),
	.B1 (n_1026),
	.B0 (ar1[7]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[7]) );
   AOI22X1 i_917 ( .Y (n_1117),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[7]),
	.A1 (dmov_inc),
	.A0 (mdr[7]) );
   OAI222XL i_915 ( .Y (n_1120),
	.C1 (n_1050),
	.C0 (n_554),
	.B1 (n_1086),
	.B0 (n_566),
	.A1 (n_1049),
	.A0 (n_548) );
   AOI31X1 i_913 ( .Y (n_1121),
	.B0 (n_922),
	.A2 (acc[8]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   AOI222X1 i_911 ( .Y (n_1124),
	.C1 (n_1015),
	.C0 (port_data_out[8]),
	.B1 (n_1026),
	.B0 (ar1[8]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[8]) );
   AOI22X1 i_909 ( .Y (n_1125),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[8]),
	.A1 (dmov_inc),
	.A0 (mdr[8]) );
   OAI222XL i_907 ( .Y (n_1128),
	.C1 (n_1050),
	.C0 (n_551),
	.B1 (n_1086),
	.B0 (n_563),
	.A1 (n_1049),
	.A0 (n_545) );
   AOI31X1 i_905 ( .Y (n_1129),
	.B0 (n_912),
	.A2 (acc[9]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   AOI222X1 i_903 ( .Y (n_1132),
	.C1 (n_1015),
	.C0 (port_data_out[9]),
	.B1 (n_1026),
	.B0 (ar1[9]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[9]) );
   AOI22X1 i_901 ( .Y (n_1133),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[9]),
	.A1 (dmov_inc),
	.A0 (mdr[9]) );
   OAI222XL i_899 ( .Y (n_1136),
	.C1 (n_1050),
	.C0 (n_548),
	.B1 (n_1086),
	.B0 (n_560),
	.A1 (n_1049),
	.A0 (n_542) );
   AOI31X1 i_897 ( .Y (n_1137),
	.B0 (n_902),
	.A2 (acc[10]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   AOI222X1 i_895 ( .Y (n_1140),
	.C1 (n_1015),
	.C0 (port_data_out[10]),
	.B1 (n_1026),
	.B0 (ar1[10]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[10]) );
   AOI22X1 i_893 ( .Y (n_1141),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[10]),
	.A1 (dmov_inc),
	.A0 (mdr[10]) );
   OAI222XL i_891 ( .Y (n_1144),
	.C1 (n_1050),
	.C0 (n_545),
	.B1 (n_1086),
	.B0 (n_557),
	.A1 (n_1049),
	.A0 (n_539) );
   AOI31X1 i_889 ( .Y (n_1145),
	.B0 (n_892),
	.A2 (acc[11]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   AOI222X1 i_887 ( .Y (n_1148),
	.C1 (n_1015),
	.C0 (port_data_out[11]),
	.B1 (n_1026),
	.B0 (ar1[11]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[11]) );
   AOI22X1 i_885 ( .Y (n_1149),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[11]),
	.A1 (dmov_inc),
	.A0 (mdr[11]) );
   NAND2X1 i_61 ( .Y (n_1152),
	.B (n_1048),
	.A (acc[28]) );
   AOI32X1 i_882 ( .Y (n_1153),
	.B1 (n_4514),
	.B0 (n_1041),
	.A2 (acc[27]),
	.A1 (n_1048),
	.A0 (n_1031) );
   OAI21XL i_883 ( .Y (n_1154),
	.B0 (n_1153),
	.A1 (n_1086),
	.A0 (n_554) );
   OAI22X1 i_880 ( .Y (n_1155),
	.B1 (n_1050),
	.B0 (n_542),
	.A1 (n_1069),
	.A0 (n_548) );
   AOI31X1 i_881 ( .Y (n_1156),
	.B0 (n_1155),
	.A2 (acc[12]),
	.A1 (FE_OFN92_n_1037),
	.A0 (n_1045) );
   AOI222X1 i_878 ( .Y (n_1159),
	.C1 (n_1015),
	.C0 (port_data_out[12]),
	.B1 (n_1026),
	.B0 (ar1[12]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[12]) );
   AOI22X1 i_876 ( .Y (n_1160),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[12]),
	.A1 (dmov_inc),
	.A0 (mdr[12]) );
   AOI32X1 i_873 ( .Y (n_1163),
	.B1 (n_4514),
	.B0 (n_1031),
	.A2 (acc[29]),
	.A1 (n_1048),
	.A0 (n_1041) );
   OAI21XL i_874 ( .Y (n_1164),
	.B0 (n_1163),
	.A1 (n_1086),
	.A0 (n_551) );
   OAI22X1 i_871 ( .Y (n_1165),
	.B1 (n_1050),
	.B0 (n_539),
	.A1 (n_1069),
	.A0 (n_545) );
   AOI31X1 i_872 ( .Y (n_1166),
	.B0 (n_1165),
	.A2 (FE_OFN92_n_1037),
	.A1 (acc[13]),
	.A0 (n_1045) );
   AOI222X1 i_869 ( .Y (n_1169),
	.C1 (n_1015),
	.C0 (port_data_out[13]),
	.B1 (n_1026),
	.B0 (ar1[13]),
	.A1 (FE_OFN94_n_1023),
	.A0 (ar0[13]) );
   AOI22X1 i_867 ( .Y (n_1170),
	.B1 (FE_OFN93_n_1035),
	.B0 (p_data_out[13]),
	.A1 (dmov_inc),
	.A0 (mdr[13]) );
   NAND2X1 i_866 ( .Y (n_1172),
	.B (n_1048),
	.A (acc[27]) );
   OAI21XL i_863 ( .Y (n_1173),
	.B0 (n_863),
	.A1 (n_1172),
	.A0 (n_452) );
   AOI31X1 i_864 ( .Y (n_1174),
	.B0 (n_1173),
	.A2 (n_1031),
	.A1 (acc[29]),
	.A0 (n_1048) );
   OAI222XL i_862 ( .Y (n_1176),
	.C1 (n_1069),
	.C0 (n_542),
	.B1 (n_4506),
	.B0 (n_1152),
	.A1 (n_1086),
	.A0 (n_548) );
   AOI222X1 i_859 ( .Y (n_1179),
	.C1 (FE_OFN94_n_1023),
	.C0 (ar0[14]),
	.B1 (n_4513),
	.B0 (acc[14]),
	.A1 (n_1026),
	.A0 (ar1[14]) );
   AOI222XL i_857 ( .Y (n_1181),
	.C1 (dmov_inc),
	.C0 (mdr[14]),
	.B1 (n_1015),
	.B0 (port_data_out[14]),
	.A1 (FE_OFN93_n_1035),
	.A0 (p_data_out[14]) );
   OAI222XL i_851 ( .Y (n_1187),
	.C1 (n_1069),
	.C0 (n_539),
	.B1 (n_1152),
	.B0 (n_452),
	.A1 (n_1086),
	.A0 (n_545) );
   NAND4BXL i_854 ( .Y (n_1188),
	.D (n_852),
	.C (n_850),
	.B (n_851),
	.AN (n_1187) );
   AOI222X1 i_848 ( .Y (n_1190),
	.C1 (FE_OFN94_n_1023),
	.C0 (ar0[15]),
	.B1 (n_4513),
	.B0 (acc[15]),
	.A1 (n_1026),
	.A0 (ar1[15]) );
   AOI222X1 i_846 ( .Y (n_1192),
	.C1 (mdr[15]),
	.C0 (dmov_inc),
	.B1 (n_1015),
	.B0 (port_data_out[15]),
	.A1 (FE_OFN93_n_1035),
	.A0 (p_data_out[15]) );
   MXI2X1 i_29 ( .Y (n_1194),
	.S0 (ir[7]),
	.B (ar[7]),
	.A (dp) );
   MXI2X1 i_578618 ( .Y (n_1195),
	.S0 (ir[7]),
	.B (ar[6]),
	.A (ir[6]) );
   MXI2X1 i_588619 ( .Y (n_1196),
	.S0 (ir[7]),
	.B (ar[5]),
	.A (ir[5]) );
   MXI2X1 i_24 ( .Y (n_1197),
	.S0 (ir[7]),
	.B (ar[4]),
	.A (ir[4]) );
   MXI2X1 i_608621 ( .Y (n_1198),
	.S0 (ir[7]),
	.B (ar_36576),
	.A (n_4524) );
   MXI2X1 i_18 ( .Y (n_1199),
	.S0 (ir[7]),
	.B (ar_26577),
	.A (n_4523) );
   MXI2X1 i_638624 ( .Y (n_1200),
	.S0 (ir[7]),
	.B (ar_06579),
	.A (n_4521) );
   MXI2X1 i_628623 ( .Y (n_1201),
	.S0 (ir[7]),
	.B (ar_16578),
	.A (n_4522) );
   NAND4X1 i_35 ( .Y (n_1204),
	.D (n_1200),
	.C (n_1201),
	.B (dmov_inc),
	.A (n_1199) );
   NOR2BX1 i_59 ( .Y (n_1205),
	.B (n_1204),
	.AN (n_1198) );
   NOR2BX1 i_17 ( .Y (n_1206),
	.B (n_1197),
	.AN (n_1205) );
   NOR2BX1 i_54 ( .Y (n_1207),
	.B (n_1196),
	.AN (n_1206) );
   NOR2BX1 i_67 ( .Y (n_1208),
	.B (n_1195),
	.AN (n_1207) );
   NAND2X1 i_55 ( .Y (n_1209),
	.B (n_1200),
	.A (dmov_inc) );
   NAND3X1 i_68 ( .Y (n_1210),
	.C (n_1201),
	.B (n_1200),
	.A (dmov_inc) );
   NOR2X1 i_56 ( .Y (n_1211),
	.B (sel_op_b[0]),
	.A (sel_op_b[2]) );
   NOR3BX1 i_2 ( .Y (n_1213),
	.C (sel_op_b[1]),
	.B (sel_op_b[0]),
	.AN (sel_op_b[2]) );
   NOR2BX1 i_841 ( .Y (n_1214),
	.B (sel_op_b[1]),
	.AN (sel_op_b[0]) );
   NOR2BX1 i_12 ( .Y (n_1215),
	.B (sel_op_b[2]),
	.AN (n_1214) );
   AOI22X1 i_840 ( .Y (n_1216),
	.B1 (n_1211),
	.B0 (mdr[15]),
	.A1 (n_1215),
	.A0 (mdr[14]) );
   NAND2X1 i_5 ( .Y (n_1217),
	.B (n_1211),
	.A (ir[11]) );
   NAND3X1 i_28 ( .Y (n_1218),
	.C (port_addrs_in[2]),
	.B (n_1211),
	.A (ir[11]) );
   AOI22X1 i_839 ( .Y (n_1219),
	.B1 (n_4511),
	.B0 (n_4496),
	.A1 (n_1215),
	.A0 (mdr[13]) );
   NOR3X1 i_3 ( .Y (n_1220),
	.C (ir[11]),
	.B (sel_op_b[0]),
	.A (sel_op_b[2]) );
   NAND2BX1 i_15 ( .Y (n_1221),
	.B (mdr[15]),
	.AN (port_addrs_in[2]) );
   OAI21XL i_52 ( .Y (n_1222),
	.B0 (n_807),
	.A1 (n_1221),
	.A0 (n_1217) );
   AOI21X1 i_838 ( .Y (n_1223),
	.B0 (n_1222),
	.A1 (n_1213),
	.A0 (p[29]) );
   AOI21X1 i_835 ( .Y (n_1226),
	.B0 (n_1222),
	.A1 (n_1213),
	.A0 (p[28]) );
   AOI22X1 i_834 ( .Y (n_1227),
	.B1 (n_1031),
	.B0 (mdr[14]),
	.A1 (n_1041),
	.A0 (mdr[15]) );
   AOI22X1 i_833 ( .Y (n_1228),
	.B1 (n_1039),
	.B0 (mdr[13]),
	.A1 (n_4508),
	.A0 (mdr[12]) );
   AOI22X1 i_832 ( .Y (n_1229),
	.B1 (n_4511),
	.B0 (n_446),
	.A1 (n_1215),
	.A0 (mdr[11]) );
   AOI21X1 i_831 ( .Y (n_1230),
	.B0 (n_1222),
	.A1 (n_1213),
	.A0 (p[27]) );
   AOI22X1 i_830 ( .Y (n_1231),
	.B1 (n_1031),
	.B0 (mdr[13]),
	.A1 (n_1041),
	.A0 (mdr[14]) );
   AOI22X1 i_829 ( .Y (n_1232),
	.B1 (n_1039),
	.B0 (mdr[12]),
	.A1 (n_4508),
	.A0 (mdr[11]) );
   AOI22X1 i_828 ( .Y (n_1233),
	.B1 (n_4511),
	.B0 (n_445),
	.A1 (n_1215),
	.A0 (mdr[10]) );
   AOI21X1 i_827 ( .Y (n_1234),
	.B0 (n_1222),
	.A1 (n_1213),
	.A0 (p[26]) );
   AOI22X1 i_826 ( .Y (n_1235),
	.B1 (n_1031),
	.B0 (mdr[12]),
	.A1 (n_1041),
	.A0 (mdr[13]) );
   AOI22X1 i_825 ( .Y (n_1236),
	.B1 (n_1039),
	.B0 (mdr[11]),
	.A1 (n_4508),
	.A0 (mdr[10]) );
   NOR2X1 i_25 ( .Y (n_1237),
	.B (n_1217),
	.A (port_addrs_in[2]) );
   AOI222X1 i_824 ( .Y (n_1239),
	.C1 (n_1215),
	.C0 (mdr[9]),
	.B1 (n_4511),
	.B0 (n_444),
	.A1 (n_4496),
	.A0 (n_1237) );
   AOI22X1 i_821 ( .Y (n_1241),
	.B1 (n_1031),
	.B0 (mdr[11]),
	.A1 (n_1041),
	.A0 (mdr[12]) );
   OAI22X1 i_818 ( .Y (n_1243),
	.B1 (n_1218),
	.B0 (n_443),
	.A1 (n_4509),
	.A0 (n_447) );
   AOI21X1 i_819 ( .Y (n_1244),
	.B0 (n_1243),
	.A1 (n_1215),
	.A0 (mdr[8]) );
   AOI22X1 i_816 ( .Y (n_1246),
	.B1 (n_1031),
	.B0 (mdr[10]),
	.A1 (n_1041),
	.A0 (mdr[11]) );
   AOI22X1 i_815 ( .Y (n_1247),
	.B1 (n_1039),
	.B0 (mdr[9]),
	.A1 (n_4508),
	.A0 (mdr[8]) );
   AOI222X1 i_814 ( .Y (n_1249),
	.C1 (n_1215),
	.C0 (mdr[7]),
	.B1 (n_4511),
	.B0 (n_442),
	.A1 (n_1237),
	.A0 (n_446) );
   AOI22X1 i_811 ( .Y (n_1251),
	.B1 (n_1031),
	.B0 (mdr[9]),
	.A1 (n_1041),
	.A0 (mdr[10]) );
   AOI22X1 i_810 ( .Y (n_1252),
	.B1 (n_1039),
	.B0 (mdr[8]),
	.A1 (n_4508),
	.A0 (mdr[7]) );
   AOI222X1 i_809 ( .Y (n_1254),
	.C1 (n_1215),
	.C0 (mdr[6]),
	.B1 (n_4511),
	.B0 (n_441),
	.A1 (n_1237),
	.A0 (n_445) );
   AOI22X1 i_806 ( .Y (n_1256),
	.B1 (n_1031),
	.B0 (mdr[8]),
	.A1 (n_1041),
	.A0 (mdr[9]) );
   AOI22X1 i_805 ( .Y (n_1257),
	.B1 (n_1039),
	.B0 (mdr[7]),
	.A1 (n_4508),
	.A0 (mdr[6]) );
   NAND2X1 i_26 ( .Y (n_1258),
	.B (n_1220),
	.A (port_addrs_in[2]) );
   AOI222X1 i_804 ( .Y (n_1260),
	.C1 (n_1237),
	.C0 (n_444),
	.B1 (n_4511),
	.B0 (n_440),
	.A1 (n_4507),
	.A0 (n_4496) );
   AOI22X1 i_801 ( .Y (n_1261),
	.B1 (n_1215),
	.B0 (mdr[5]),
	.A1 (n_1213),
	.A0 (p[21]) );
   AOI22X1 i_800 ( .Y (n_1263),
	.B1 (n_1031),
	.B0 (mdr[7]),
	.A1 (n_1041),
	.A0 (mdr[8]) );
   AOI22X1 i_799 ( .Y (n_1264),
	.B1 (n_1039),
	.B0 (mdr[6]),
	.A1 (n_4508),
	.A0 (mdr[5]) );
   OAI222XL i_798 ( .Y (n_1266),
	.C1 (n_4509),
	.C0 (n_443),
	.B1 (n_4498),
	.B0 (n_1218),
	.A1 (n_1258),
	.A0 (n_447) );
   AOI22X1 i_795 ( .Y (n_1267),
	.B1 (n_1215),
	.B0 (mdr[4]),
	.A1 (n_1213),
	.A0 (p[20]) );
   AOI22X1 i_794 ( .Y (n_1269),
	.B1 (n_1031),
	.B0 (mdr[6]),
	.A1 (n_1041),
	.A0 (mdr[7]) );
   AOI22X1 i_793 ( .Y (n_1270),
	.B1 (n_1039),
	.B0 (mdr[5]),
	.A1 (n_4508),
	.A0 (mdr[4]) );
   AOI211X1 i_792 ( .Y (n_1272),
	.C0 (n_757),
	.B0 (n_758),
	.A1 (n_1237),
	.A0 (n_442) );
   AOI22X1 i_789 ( .Y (n_1273),
	.B1 (n_1215),
	.B0 (mdr[3]),
	.A1 (n_1213),
	.A0 (p[19]) );
   AOI22X1 i_788 ( .Y (n_1275),
	.B1 (n_1031),
	.B0 (mdr[5]),
	.A1 (n_1041),
	.A0 (mdr[6]) );
   AOI22X1 i_787 ( .Y (n_1276),
	.B1 (n_1039),
	.B0 (mdr[4]),
	.A1 (n_4508),
	.A0 (mdr[3]) );
   AOI222X1 i_786 ( .Y (n_1278),
	.C1 (n_1237),
	.C0 (n_441),
	.B1 (n_4511),
	.B0 (n_437),
	.A1 (n_4507),
	.A0 (n_445) );
   AOI22X1 i_783 ( .Y (n_1279),
	.B1 (n_1215),
	.B0 (mdr[2]),
	.A1 (n_1213),
	.A0 (p[18]) );
   AOI22X1 i_782 ( .Y (n_1281),
	.B1 (n_1031),
	.B0 (mdr[4]),
	.A1 (n_1041),
	.A0 (mdr[5]) );
   AOI22X1 i_781 ( .Y (n_1282),
	.B1 (n_1039),
	.B0 (mdr[3]),
	.A1 (n_4508),
	.A0 (mdr[2]) );
   NAND2BX1 i_27 ( .Y (n_1283),
	.B (n_1220),
	.AN (port_addrs_in[2]) );
   OAI222XL i_780 ( .Y (n_1285),
	.C1 (n_4497),
	.C0 (n_1258),
	.B1 (n_1218),
	.B0 (n_4499),
	.A1 (n_449),
	.A0 (n_1283) );
   AOI222X1 i_778 ( .Y (n_1287),
	.C1 (n_1213),
	.C0 (p[17]),
	.B1 (n_1237),
	.B0 (n_440),
	.A1 (n_1215),
	.A0 (mdr[1]) );
   AOI22X1 i_776 ( .Y (n_1288),
	.B1 (n_1031),
	.B0 (mdr[3]),
	.A1 (n_1041),
	.A0 (mdr[4]) );
   AOI22X1 i_775 ( .Y (n_1289),
	.B1 (n_1039),
	.B0 (mdr[2]),
	.A1 (n_4508),
	.A0 (mdr[1]) );
   OAI222XL i_774 ( .Y (n_1291),
	.C1 (n_443),
	.C0 (n_1258),
	.B1 (n_4500),
	.B0 (n_1218),
	.A1 (n_1283),
	.A0 (n_447) );
   AOI222X1 i_772 ( .Y (n_1293),
	.C1 (n_1213),
	.C0 (p[16]),
	.B1 (n_439),
	.B0 (n_1237),
	.A1 (n_1215),
	.A0 (mdr[0]) );
   AOI22X1 i_770 ( .Y (n_1294),
	.B1 (n_1031),
	.B0 (mdr[2]),
	.A1 (n_1041),
	.A0 (mdr[3]) );
   AOI22X1 i_767 ( .Y (n_1295),
	.B1 (n_430),
	.B0 (n_4511),
	.A1 (n_4505),
	.A0 (n_446) );
   AOI22X1 i_766 ( .Y (n_1296),
	.B1 (n_4507),
	.B0 (n_442),
	.A1 (n_1237),
	.A0 (n_438) );
   NAND2X1 i_11 ( .Y (n_1298),
	.B (n_1214),
	.A (sel_op_b[2]) );
   NOR2BX1 i_10 ( .Y (n_1299),
	.B (n_1211),
	.AN (sel_op_b[1]) );
   AOI22X1 i_764 ( .Y (n_1300),
	.B1 (n_1299),
	.B0 (mdr[15]),
	.A1 (n_1213),
	.A0 (p[15]) );
   AOI22X1 i_761 ( .Y (n_1303),
	.B1 (n_4502),
	.B0 (n_4511),
	.A1 (n_4505),
	.A0 (n_445) );
   AOI22X1 i_760 ( .Y (n_1304),
	.B1 (n_4507),
	.B0 (n_441),
	.A1 (n_1237),
	.A0 (n_437) );
   AOI22X1 i_758 ( .Y (n_1306),
	.B1 (n_1299),
	.B0 (mdr[14]),
	.A1 (n_1213),
	.A0 (p[14]) );
   NOR2X1 i_64 ( .Y (n_1308),
	.B (port_addrs_in[1]),
	.A (n_432) );
   AOI22X1 i_756 ( .Y (n_1309),
	.B1 (n_4511),
	.B0 (n_1308),
	.A1 (n_4505),
	.A0 (n_444) );
   AOI22X1 i_755 ( .Y (n_1310),
	.B1 (n_4507),
	.B0 (n_440),
	.A1 (n_436),
	.A0 (n_1237) );
   AOI22X1 i_753 ( .Y (n_1312),
	.B1 (n_1299),
	.B0 (mdr[13]),
	.A1 (n_1213),
	.A0 (p[13]) );
   NAND2X1 i_34 ( .Y (n_1314),
	.B (n_1041),
	.A (mdr[0]) );
   AOI2BB1X1 i_751 ( .Y (n_1315),
	.B0 (n_701),
	.A1N (n_1283),
	.A0N (n_443) );
   AOI22X1 i_750 ( .Y (n_1316),
	.B1 (n_4507),
	.B0 (n_439),
	.A1 (n_1237),
	.A0 (n_435) );
   AOI22X1 i_748 ( .Y (n_1318),
	.B1 (n_1299),
	.B0 (mdr[12]),
	.A1 (n_1213),
	.A0 (p[12]) );
   AOI22X1 i_746 ( .Y (n_1320),
	.B1 (n_4505),
	.B0 (n_442),
	.A1 (n_4507),
	.A0 (n_438) );
   AOI222X1 i_745 ( .Y (n_1323),
	.C1 (n_1213),
	.C0 (p[11]),
	.B1 (n_4504),
	.B0 (ir[11]),
	.A1 (n_1299),
	.A0 (mdr[11]) );
   AOI22X1 i_742 ( .Y (n_1324),
	.B1 (n_4505),
	.B0 (n_441),
	.A1 (n_4507),
	.A0 (n_437) );
   AOI222X1 i_741 ( .Y (n_1327),
	.C1 (n_1213),
	.C0 (p[10]),
	.B1 (n_4504),
	.B0 (port_addrs_in[2]),
	.A1 (n_1299),
	.A0 (mdr[10]) );
   AOI22X1 i_738 ( .Y (n_1328),
	.B1 (n_1237),
	.B0 (n_1308),
	.A1 (n_4505),
	.A0 (n_440) );
   AOI222X1 i_737 ( .Y (n_1331),
	.C1 (n_1213),
	.C0 (p[9]),
	.B1 (n_4504),
	.B0 (port_addrs_in[1]),
	.A1 (n_1299),
	.A0 (mdr[9]) );
   AOI22X1 i_734 ( .Y (n_1332),
	.B1 (n_4505),
	.B0 (n_439),
	.A1 (n_435),
	.A0 (n_4507) );
   AOI222X1 i_733 ( .Y (n_1335),
	.C1 (n_1213),
	.C0 (p[8]),
	.B1 (n_4504),
	.B0 (port_addrs_in[0]),
	.A1 (n_1299),
	.A0 (mdr[8]) );
   AOI22X1 i_730 ( .Y (n_1336),
	.B1 (n_4505),
	.B0 (n_438),
	.A1 (n_4507),
	.A0 (n_430) );
   AOI22X1 i_729 ( .Y (n_1338),
	.B1 (n_1299),
	.B0 (mdr[7]),
	.A1 (n_1213),
	.A0 (p[7]) );
   AOI22X1 i_727 ( .Y (n_1339),
	.B1 (n_4505),
	.B0 (n_437),
	.A1 (n_4507),
	.A0 (n_4502) );
   AOI22X1 i_726 ( .Y (n_1341),
	.B1 (n_1299),
	.B0 (mdr[6]),
	.A1 (n_1213),
	.A0 (p[6]) );
   OAI21XL i_724 ( .Y (n_1342),
	.B0 (n_660),
	.A1 (n_1283),
	.A0 (n_4499) );
   AOI31X1 i_725 ( .Y (n_1343),
	.B0 (n_1342),
	.A2 (n_1214),
	.A1 (ir[5]),
	.A0 (sel_op_b[2]) );
   AOI22X1 i_723 ( .Y (n_1344),
	.B1 (n_1299),
	.B0 (mdr[5]),
	.A1 (n_1213),
	.A0 (p[5]) );
   AOI32X1 i_721 ( .Y (n_1345),
	.B1 (n_4505),
	.B0 (n_435),
	.A2 (n_4507),
	.A1 (n_1041),
	.A0 (mdr[0]) );
   AOI22X1 i_720 ( .Y (n_1347),
	.B1 (n_1299),
	.B0 (mdr[4]),
	.A1 (n_1213),
	.A0 (p[4]) );
   AOI22X1 i_718 ( .Y (n_1349),
	.B1 (n_1299),
	.B0 (mdr[3]),
	.A1 (n_1213),
	.A0 (p[3]) );
   AOI22X1 i_716 ( .Y (n_1351),
	.B1 (n_1299),
	.B0 (mdr[2]),
	.A1 (n_1213),
	.A0 (p[2]) );
   AOI32X1 i_715 ( .Y (n_1352),
	.B1 (n_4505),
	.B0 (n_1308),
	.A2 (ir[1]),
	.A1 (n_1214),
	.A0 (sel_op_b[2]) );
   AOI22X1 i_714 ( .Y (n_1353),
	.B1 (n_1299),
	.B0 (mdr[1]),
	.A1 (n_1213),
	.A0 (p[1]) );
   AOI22X1 i_712 ( .Y (n_1355),
	.B1 (n_1299),
	.B0 (mdr[0]),
	.A1 (n_1213),
	.A0 (p[0]) );
   NOR3BX1 i_1 ( .Y (n_1357),
	.C (sel_op_a[2]),
	.B (sel_op_a[1]),
	.AN (sel_op_a[0]) );
   NAND2X1 i_710 ( .Y (n_1358),
	.B (sel_op_a[0]),
	.A (sel_op_a[1]) );
   NOR2X1 i_8 ( .Y (n_1359),
	.B (sel_op_a[2]),
	.A (n_1358) );
   AOI22X1 i_709 ( .Y (n_1360),
	.B1 (n_1359),
	.B0 (top[15]),
	.A1 (n_1357),
	.A0 (acc[15]) );
   AOI22X1 i_708 ( .Y (n_1361),
	.B1 (n_1359),
	.B0 (top[14]),
	.A1 (n_1357),
	.A0 (acc[14]) );
   AOI22X1 i_707 ( .Y (n_1362),
	.B1 (n_1359),
	.B0 (top[13]),
	.A1 (n_1357),
	.A0 (acc[13]) );
   AOI22X1 i_706 ( .Y (n_1363),
	.B1 (n_1359),
	.B0 (top[12]),
	.A1 (n_1357),
	.A0 (acc[12]) );
   AOI22X1 i_705 ( .Y (n_1364),
	.B1 (n_1359),
	.B0 (top[11]),
	.A1 (n_1357),
	.A0 (acc[11]) );
   AOI22X1 i_704 ( .Y (n_1365),
	.B1 (n_1359),
	.B0 (top[10]),
	.A1 (n_1357),
	.A0 (acc[10]) );
   AOI22X1 i_703 ( .Y (n_1366),
	.B1 (n_1359),
	.B0 (top[9]),
	.A1 (n_1357),
	.A0 (acc[9]) );
   AOI22X1 i_702 ( .Y (n_1367),
	.B1 (n_1359),
	.B0 (top[8]),
	.A1 (n_1357),
	.A0 (acc[8]) );
   NOR2X1 i_14 ( .Y (n_1368),
	.B (n_4520),
	.A (n_1358) );
   AOI22X1 i_700 ( .Y (n_1369),
	.B1 (n_1368),
	.B0 (ir[7]),
	.A1 (n_1359),
	.A0 (top[7]) );
   AOI22X1 i_699 ( .Y (n_1370),
	.B1 (n_1357),
	.B0 (acc[7]),
	.A1 (n_410),
	.A0 (mdr[7]) );
   AOI22X1 i_698 ( .Y (n_1371),
	.B1 (n_1368),
	.B0 (ir[6]),
	.A1 (n_1359),
	.A0 (top[6]) );
   AOI22X1 i_697 ( .Y (n_1372),
	.B1 (n_1357),
	.B0 (acc[6]),
	.A1 (n_410),
	.A0 (mdr[6]) );
   AOI22X1 i_696 ( .Y (n_1373),
	.B1 (n_1368),
	.B0 (ir[5]),
	.A1 (n_1359),
	.A0 (top[5]) );
   AOI22X1 i_695 ( .Y (n_1374),
	.B1 (n_1357),
	.B0 (acc[5]),
	.A1 (n_410),
	.A0 (mdr[5]) );
   AOI22X1 i_694 ( .Y (n_1375),
	.B1 (n_1368),
	.B0 (ir[4]),
	.A1 (n_1359),
	.A0 (top[4]) );
   AOI22X1 i_693 ( .Y (n_1376),
	.B1 (n_1357),
	.B0 (acc[4]),
	.A1 (n_410),
	.A0 (mdr[4]) );
   AOI22X1 i_691 ( .Y (n_1378),
	.B1 (n_1357),
	.B0 (acc[3]),
	.A1 (n_410),
	.A0 (mdr[3]) );
   AOI22X1 i_689 ( .Y (n_1380),
	.B1 (n_1357),
	.B0 (acc[2]),
	.A1 (n_410),
	.A0 (mdr[2]) );
   AOI22X1 i_688 ( .Y (n_1381),
	.B1 (n_1368),
	.B0 (ir[1]),
	.A1 (n_1359),
	.A0 (top[1]) );
   AOI22X1 i_687 ( .Y (n_1382),
	.B1 (acc[1]),
	.B0 (n_1357),
	.A1 (n_410),
	.A0 (mdr[1]) );
   AOI22X1 i_685 ( .Y (n_1384),
	.B1 (acc[0]),
	.B0 (n_1357),
	.A1 (n_410),
	.A0 (mdr[0]) );
   OR2X1 i_5354 ( .Y (go_prog),
	.B (dec_go_prog),
	.A (enc_go_prog) );
   OR2X1 i_5356 ( .Y (go_port),
	.B (dec_go_port),
	.A (enc_go_port) );
   OR2X1 i_5357 ( .Y (go_data),
	.B (dec_go_data),
	.A (enc_go_data) );
   OR2X1 i_5358 ( .Y (read_data),
	.B (dec_read_data),
	.A (enc_read_data) );
   OR2X1 i_5366 ( .Y (read_prog),
	.B (dec_read_prog),
	.A (enc_read_prog) );
   OR2X1 i_5369 ( .Y (read_port),
	.B (dec_read_port),
	.A (enc_read_port) );
   NAND4BXL i_5427 ( .Y (data_in[0]),
	.D (n_1044),
	.C (n_1055),
	.B (n_1056),
	.AN (n_1052) );
   NAND4BXL i_5434 ( .Y (data_in[1]),
	.D (n_1059),
	.C (n_1064),
	.B (n_1065),
	.AN (n_1061) );
   NAND4BXL i_5441 ( .Y (data_in[2]),
	.D (n_1071),
	.C (n_1074),
	.B (n_1075),
	.AN (n_1068) );
   NAND4BXL i_5448 ( .Y (data_in[3]),
	.D (n_1080),
	.C (n_1083),
	.B (n_1084),
	.AN (n_1078) );
   NAND4BXL i_5455 ( .Y (data_in[4]),
	.D (n_1089),
	.C (n_1092),
	.B (n_1093),
	.AN (n_1088) );
   NAND4BXL i_5462 ( .Y (data_in[5]),
	.D (n_1097),
	.C (n_1100),
	.B (n_1101),
	.AN (n_1096) );
   NAND4BXL i_5469 ( .Y (data_in[6]),
	.D (n_1105),
	.C (n_1108),
	.B (n_1109),
	.AN (n_1104) );
   NAND4BXL i_5476 ( .Y (data_in[7]),
	.D (n_1113),
	.C (n_1116),
	.B (n_1117),
	.AN (n_1112) );
   NAND4BXL i_5483 ( .Y (data_in[8]),
	.D (n_1121),
	.C (n_1124),
	.B (n_1125),
	.AN (n_1120) );
   NAND4BXL i_5490 ( .Y (data_in[9]),
	.D (n_1129),
	.C (n_1132),
	.B (n_1133),
	.AN (n_1128) );
   NAND4BXL i_5497 ( .Y (data_in[10]),
	.D (n_1137),
	.C (n_1140),
	.B (n_1141),
	.AN (n_1136) );
   NAND4BXL i_5504 ( .Y (data_in[11]),
	.D (n_1145),
	.C (n_1148),
	.B (n_1149),
	.AN (n_1144) );
   NAND4BXL i_5511 ( .Y (data_in[12]),
	.D (n_1156),
	.C (n_1159),
	.B (n_1160),
	.AN (n_1154) );
   NAND4BXL i_5518 ( .Y (data_in[13]),
	.D (n_1166),
	.C (n_1169),
	.B (n_1170),
	.AN (n_1164) );
   NAND4BXL i_5525 ( .Y (data_in[14]),
	.D (n_1174),
	.C (n_1179),
	.B (n_1181),
	.AN (n_1176) );
   NAND3BX1 i_5532 ( .Y (data_in[15]),
	.C (n_1190),
	.B (n_1192),
	.AN (n_1188) );
   MX2X1 i_248287 ( .Y (ar[15]),
	.S0 (arp),
	.B (ar1[15]),
	.A (ar0[15]) );
   MX2X1 i_258288 ( .Y (ar[14]),
	.S0 (arp),
	.B (ar1[14]),
	.A (ar0[14]) );
   MX2X1 i_268289 ( .Y (ar[13]),
	.S0 (arp),
	.B (ar1[13]),
	.A (ar0[13]) );
   MX2X1 i_278290 ( .Y (ar[12]),
	.S0 (arp),
	.B (ar1[12]),
	.A (ar0[12]) );
   MX2X1 i_288291 ( .Y (ar[11]),
	.S0 (arp),
	.B (ar1[11]),
	.A (ar0[11]) );
   MX2X1 i_298292 ( .Y (ar[10]),
	.S0 (arp),
	.B (ar1[10]),
	.A (ar0[10]) );
   MX2X1 i_308293 ( .Y (ar[9]),
	.S0 (arp),
	.B (ar1[9]),
	.A (ar0[9]) );
   MX2X1 i_318294 ( .Y (ar[8]),
	.S0 (arp),
	.B (ar1[8]),
	.A (ar0[8]) );
   MX2X1 i_328295 ( .Y (ar[7]),
	.S0 (arp),
	.B (ar1[7]),
	.A (ar0[7]) );
   MX2X1 i_338296 ( .Y (ar[6]),
	.S0 (arp),
	.B (ar1[6]),
	.A (ar0[6]) );
   MX2X1 i_348297 ( .Y (ar[5]),
	.S0 (arp),
	.B (ar1[5]),
	.A (ar0[5]) );
   MX2X1 i_358298 ( .Y (ar[4]),
	.S0 (arp),
	.B (ar1[4]),
	.A (ar0[4]) );
   MXI2X1 i_368299 ( .Y (ar_36576),
	.S0 (arp),
	.B (ar1[3]),
	.A (ar0[3]) );
   MXI2X1 i_378300 ( .Y (ar_26577),
	.S0 (arp),
	.B (ar1[2]),
	.A (ar0[2]) );
   MXI2X1 i_388301 ( .Y (ar_16578),
	.S0 (arp),
	.B (ar1[1]),
	.A (ar0[1]) );
   MXI2X1 i_398302 ( .Y (ar_06579),
	.S0 (arp),
	.B (ar1[0]),
	.A (ar0[0]) );
   OAI21XL i_568625 ( .Y (addrs_in[7]),
	.B0 (n_489),
	.A1 (n_1194),
	.A0 (n_1208) );
   OAI21XL i_578626 ( .Y (addrs_in[6]),
	.B0 (n_487),
	.A1 (n_1195),
	.A0 (n_1207) );
   OAI21XL i_588627 ( .Y (addrs_in[5]),
	.B0 (n_485),
	.A1 (n_1196),
	.A0 (n_1206) );
   OAI21XL i_598628 ( .Y (addrs_in[4]),
	.B0 (n_483),
	.A1 (n_1197),
	.A0 (n_1205) );
   OAI21XL i_608629 ( .Y (addrs_in[3]),
	.B0 (n_482),
	.A1 (n_1198),
	.A0 (n_1204) );
   OAI21XL i_618630 ( .Y (addrs_in[2]),
	.B0 (n_480),
	.A1 (n_1199),
	.A0 (n_1210) );
   OAI21XL i_628631 ( .Y (addrs_in[1]),
	.B0 (n_478),
	.A1 (n_1201),
	.A0 (n_1209) );
   XOR2X1 i_638632 ( .Y (addrs_in[0]),
	.B (dmov_inc),
	.A (n_1200) );
   MX2X1 i_582 ( .Y (p_addrs_in[7]),
	.S0 (pc_acc),
	.B (acc[7]),
	.A (pc[7]) );
   MX2X1 i_583 ( .Y (p_addrs_in[6]),
	.S0 (pc_acc),
	.B (acc[6]),
	.A (pc[6]) );
   MX2X1 i_584 ( .Y (p_addrs_in[5]),
	.S0 (pc_acc),
	.B (acc[5]),
	.A (pc[5]) );
   MX2X1 i_585 ( .Y (p_addrs_in[4]),
	.S0 (pc_acc),
	.B (acc[4]),
	.A (pc[4]) );
   MX2X1 i_586 ( .Y (p_addrs_in[3]),
	.S0 (pc_acc),
	.B (acc[3]),
	.A (pc[3]) );
   MX2X1 i_587 ( .Y (p_addrs_in[2]),
	.S0 (pc_acc),
	.B (acc[2]),
	.A (pc[2]) );
   MX2X1 i_588 ( .Y (p_addrs_in[1]),
	.S0 (pc_acc),
	.B (acc[1]),
	.A (pc[1]) );
   MX2X1 i_589 ( .Y (p_addrs_in[0]),
	.S0 (pc_acc),
	.B (acc[0]),
	.A (pc[0]) );
   AOI22X1 i_517 ( .Y (opb_316580),
	.B1 (n_456),
	.B0 (mdr[15]),
	.A1 (n_1213),
	.A0 (p[31]) );
   OAI2BB1X1 i_518 ( .Y (opb[30]),
	.B0 (n_1216),
	.A1N (n_1213),
	.A0N (p[30]) );
   NAND2X1 i_519 ( .Y (opb[29]),
	.B (n_1219),
	.A (n_1223) );
   OAI211X1 i_520 ( .Y (opb[28]),
	.C0 (n_1226),
	.B0 (n_832),
	.A1 (n_1218),
	.A0 (n_447) );
   NAND2X1 i_521 ( .Y (opb[27]),
	.B (n_1229),
	.A (n_1230) );
   NAND2X1 i_522 ( .Y (opb[26]),
	.B (n_1233),
	.A (n_1234) );
   NAND3X1 i_523 ( .Y (opb[25]),
	.C (n_1239),
	.B (n_807),
	.A (n_808) );
   NAND3X1 i_524 ( .Y (opb[24]),
	.C (n_1244),
	.B (n_799),
	.A (n_807) );
   NAND3X1 i_525 ( .Y (opb[23]),
	.C (n_1249),
	.B (n_791),
	.A (n_807) );
   NAND3X1 i_526 ( .Y (opb[22]),
	.C (n_1254),
	.B (n_783),
	.A (n_807) );
   NAND3X1 i_527 ( .Y (opb[21]),
	.C (n_1260),
	.B (n_1261),
	.A (n_775) );
   NAND3X1 i_528 ( .Y (opb[20]),
	.C (n_4512),
	.B (n_1267),
	.A (n_775) );
   NAND3X1 i_529 ( .Y (opb[19]),
	.C (n_1272),
	.B (n_1273),
	.A (n_775) );
   NAND3X1 i_530 ( .Y (opb[18]),
	.C (n_1278),
	.B (n_1279),
	.A (n_775) );
   NAND2BX1 i_531 ( .Y (opb[17]),
	.B (n_1287),
	.AN (n_1285) );
   NAND2BX1 i_532 ( .Y (opb[16]),
	.B (n_1293),
	.AN (n_1291) );
   NAND4X1 i_533 ( .Y (opb[15]),
	.D (n_1295),
	.C (n_1296),
	.B (n_1300),
	.A (n_719) );
   NAND4X1 i_534 ( .Y (opb[14]),
	.D (n_1303),
	.C (n_1304),
	.B (n_1306),
	.A (n_719) );
   NAND4X1 i_535 ( .Y (opb[13]),
	.D (n_1309),
	.C (n_1310),
	.B (n_1312),
	.A (n_719) );
   NAND4X1 i_536 ( .Y (opb[12]),
	.D (n_1315),
	.C (n_1316),
	.B (n_1318),
	.A (n_719) );
   OAI211X1 i_537 ( .Y (opb[11]),
	.C0 (n_1323),
	.B0 (n_1320),
	.A1 (n_4509),
	.A0 (n_4501) );
   OAI211X1 i_538 ( .Y (opb[10]),
	.C0 (n_1327),
	.B0 (n_1324),
	.A1 (n_4509),
	.A0 (n_428) );
   OAI211X1 i_539 ( .Y (opb[9]),
	.C0 (n_1331),
	.B0 (n_1328),
	.A1 (n_4499),
	.A0 (n_1258) );
   OAI211X1 i_540 ( .Y (opb[8]),
	.C0 (n_1335),
	.B0 (n_1332),
	.A1 (n_4509),
	.A0 (n_1314) );
   NAND3X1 i_541 ( .Y (opb[7]),
	.C (n_1336),
	.B (n_1338),
	.A (n_672) );
   NAND3X1 i_542 ( .Y (opb[6]),
	.C (n_1339),
	.B (n_1341),
	.A (n_667) );
   NAND2X1 i_543 ( .Y (opb[5]),
	.B (n_1343),
	.A (n_1344) );
   NAND3X1 i_544 ( .Y (opb[4]),
	.C (n_1345),
	.B (n_1347),
	.A (n_657) );
   OAI221XL i_545 ( .Y (opb[3]),
	.C0 (n_1349),
	.B1 (n_1283),
	.B0 (n_4501),
	.A1 (n_4524),
	.A0 (n_1298) );
   OAI221XL i_546 ( .Y (opb[2]),
	.C0 (n_1351),
	.B1 (n_1283),
	.B0 (n_428),
	.A1 (n_4523),
	.A0 (n_1298) );
   NAND2X1 i_547 ( .Y (opb[1]),
	.B (n_1352),
	.A (n_1353) );
   OAI221XL i_548 ( .Y (opb[0]),
	.C0 (n_1355),
	.B1 (n_1283),
	.B0 (n_1314),
	.A1 (n_4521),
	.A0 (n_1298) );
   OAI2BB1X1 i_5178960 ( .Y (opa[31]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[31]) );
   OAI2BB1X1 i_5188961 ( .Y (opa[30]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[30]) );
   OAI2BB1X1 i_5198962 ( .Y (opa[29]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[29]) );
   OAI2BB1X1 i_5208963 ( .Y (opa[28]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[28]) );
   OAI2BB1X1 i_5218964 ( .Y (opa[27]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[27]) );
   OAI2BB1X1 i_5228965 ( .Y (opa[26]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[26]) );
   OAI2BB1X1 i_5238966 ( .Y (opa[25]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[25]) );
   OAI2BB1X1 i_5248967 ( .Y (opa[24]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[24]) );
   OAI2BB1X1 i_5258968 ( .Y (opa[23]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[23]) );
   OAI2BB1X1 i_5268969 ( .Y (opa[22]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[22]) );
   OAI2BB1X1 i_5278970 ( .Y (opa[21]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[21]) );
   OAI2BB1X1 i_5288971 ( .Y (opa[20]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[20]) );
   OAI2BB1X1 i_5298972 ( .Y (opa[19]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[19]) );
   OAI2BB1X1 i_5308973 ( .Y (opa[18]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[18]) );
   OAI2BB1X1 i_5318974 ( .Y (opa[17]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[17]) );
   OAI2BB1X1 i_5328975 ( .Y (opa[16]),
	.B0 (n_402),
	.A1N (n_1357),
	.A0N (acc[16]) );
   NAND2X1 i_5338976 ( .Y (opa[15]),
	.B (n_1360),
	.A (n_402) );
   OAI2BB1X1 i_5348977 ( .Y (opa[14]),
	.B0 (n_1361),
	.A1N (n_410),
	.A0N (mdr[14]) );
   OAI2BB1X1 i_5358978 ( .Y (opa[13]),
	.B0 (n_1362),
	.A1N (n_410),
	.A0N (mdr[13]) );
   OAI2BB1X1 i_5368979 ( .Y (opa[12]),
	.B0 (n_1363),
	.A1N (n_410),
	.A0N (mdr[12]) );
   OAI2BB1X1 i_5378980 ( .Y (opa[11]),
	.B0 (n_1364),
	.A1N (n_410),
	.A0N (mdr[11]) );
   OAI2BB1X1 i_5388981 ( .Y (opa[10]),
	.B0 (n_1365),
	.A1N (n_410),
	.A0N (mdr[10]) );
   OAI2BB1X1 i_5398982 ( .Y (opa[9]),
	.B0 (n_1366),
	.A1N (n_410),
	.A0N (mdr[9]) );
   OAI2BB1X1 i_5408983 ( .Y (opa[8]),
	.B0 (n_1367),
	.A1N (n_410),
	.A0N (mdr[8]) );
   NAND2X1 i_5418984 ( .Y (opa[7]),
	.B (n_1369),
	.A (n_1370) );
   NAND2X1 i_5428985 ( .Y (opa[6]),
	.B (n_1371),
	.A (n_1372) );
   NAND2X1 i_5438986 ( .Y (opa[5]),
	.B (n_1373),
	.A (n_1374) );
   NAND2X1 i_5448987 ( .Y (opa[4]),
	.B (n_1375),
	.A (n_1376) );
   OAI211X1 i_5458988 ( .Y (opa[3]),
	.C0 (n_1378),
	.B0 (n_604),
	.A1 (n_4524),
	.A0 (n_4503) );
   OAI211X1 i_5468989 ( .Y (opa[2]),
	.C0 (n_1380),
	.B0 (n_600),
	.A1 (n_4523),
	.A0 (n_4503) );
   NAND2X1 i_5478990 ( .Y (opa[1]),
	.B (n_1381),
	.A (n_1382) );
   OAI211X1 i_5488991 ( .Y (opa[0]),
	.C0 (n_1384),
	.B0 (n_592),
	.A1 (n_4521),
	.A0 (n_4503) );
   INVX1 i_6102 ( .Y (n_4496),
	.A (n_449) );
   INVX1 i_6103 ( .Y (n_4497),
	.A (n_444) );
   INVX1 i_6104 ( .Y (n_4498),
	.A (n_439) );
   INVX1 i_6105 ( .Y (n_4499),
	.A (n_436) );
   INVX1 i_6106 ( .Y (n_4500),
	.A (n_435) );
   INVX1 i_6107 ( .Y (n_4501),
	.A (n_430) );
   INVX1 i_6108 ( .Y (n_4502),
	.A (n_428) );
   INVX1 i_6109 ( .Y (n_4503),
	.A (n_1368) );
   INVX1 i_6110 ( .Y (n_4504),
	.A (n_1298) );
   INVX1 i_6111 ( .Y (n_4505),
	.A (n_1283) );
   INVX1 i_6112 ( .Y (n_4506),
	.A (n_1039) );
   INVX1 i_6113 ( .Y (n_4507),
	.A (n_1258) );
   INVX1 i_6114 ( .Y (n_4508),
	.A (n_452) );
   INVX1 i_6115 ( .Y (n_4509),
	.A (n_1237) );
   INVX1 i_6116 ( .Y (n_4510),
	.A (n_1241) );
   INVX1 i_6117 ( .Y (n_4511),
	.A (n_1218) );
   INVX1 i_6118 ( .Y (n_4512),
	.A (n_1266) );
   INVX1 i_6119 ( .Y (n_4513),
	.A (n_1046) );
   INVX1 i_6120 ( .Y (n_4514),
	.A (n_1152) );
   INVX1 i_6121 ( .Y (opb[31]),
	.A (opb_316580) );
   INVX1 i_6122 ( .Y (ar[0]),
	.A (ar_06579) );
   INVX1 i_6123 ( .Y (ar[1]),
	.A (ar_16578) );
   INVX1 i_6124 ( .Y (ar[2]),
	.A (ar_26577) );
   INVX1 i_6125 ( .Y (ar[3]),
	.A (ar_36576) );
   INVX1 i_6126 ( .Y (n_4520),
	.A (sel_op_a[2]) );
   INVX1 i_6127 ( .Y (n_4521),
	.A (ir[0]) );
   INVX1 i_6128 ( .Y (n_4522),
	.A (ir[1]) );
   INVX1 i_6129 ( .Y (n_4523),
	.A (ir[2]) );
   INVX1 i_6130 ( .Y (n_4524),
	.A (ir[3]) );
   INVX1 i_6131 ( .Y (n_4525),
	.A (port_addrs_in[1]) );
   INVX1 i_6132 ( .Y (n_4526),
	.A (acc[0]) );
   INVX1 i_6133 ( .Y (n_4527),
	.A (acc[1]) );
   BUFX1 FE_OFC94_n_1023 ( .Y (FE_OFN94_n_1023),
	.A (n_1023) );
   BUFX1 FE_OFC93_n_1035 ( .Y (FE_OFN93_n_1035),
	.A (n_1035) );
   BUFX1 FE_OFC92_n_1037 ( .Y (FE_OFN92_n_1037),
	.A (n_1037) );
endmodule

module tdsp_core_mach (
	samp_bio,
	samp_int,
	phi_1,
	phi_2,
	phi_3,
	phi_4,
	phi_5,
	phi_6,
	reset,
	clk,
	bus_request,
	bus_grant,
	bio,
	int,
	scan_en,
	BG_scan_in,
	BG_scan_out );
   output samp_bio;
   output samp_int;
   output phi_1;
   output phi_2;
   output phi_3;
   output phi_4;
   output phi_5;
   output phi_6;
   input reset;
   input clk;
   input bus_request;
   input bus_grant;
   input bio;
   input int;
   input scan_en;
   input BG_scan_in;
   output BG_scan_out;

   // Internal wires
   wire [2:0] tdsp_state;
   wire n_102;
   wire n_47;
   wire n_27;
   wire n_45;
   wire n_72;
   wire n_22;
   wire n_23;
   wire n_24;
   wire n_35;
   wire n_2818;
   wire n_37;
   wire n_34;
   wire n_28;
   wire n_31;
   wire n_49;
   wire n_33;
   wire n_36;
   wire n_40;
   wire n_57;
   wire n_117;
   wire n_42;
   wire n_48;
   wire n_2820;
   wire n_2782;
   wire n_2822;
   wire n_2784;
   wire n_2788;
   wire n_2821;
   wire n_2790;
   wire n_2794;
   wire n_2819;
   wire n_2797;
   wire n_2800;
   wire n_2803;
   wire n_2806;
   wire n_2812;
   wire n_2815;

   CLKBUFXL i_10014 ( .Y (phi_6),
	.A (BG_scan_out) );
   NAND2X1 i_12 ( .Y (n_27),
	.B (n_47),
	.A (n_102) );
   NAND4BXL i_122 ( .Y (n_24),
	.D (n_23),
	.C (n_22),
	.B (n_72),
	.AN (n_45) );
   NAND2X1 i_14 ( .Y (n_23),
	.B (n_2818),
	.A (n_35) );
   AOI32X1 i_228675 ( .Y (n_22),
	.B1 (n_37),
	.B0 (n_35),
	.A2 (tdsp_state[0]),
	.A1 (tdsp_state[1]),
	.A0 (tdsp_state[2]) );
   NAND3X1 i_41 ( .Y (n_28),
	.C (n_34),
	.B (n_72),
	.A (n_23) );
   AOI21X1 i_5 ( .Y (n_31),
	.B0 (tdsp_state[0]),
	.A1 (bus_grant),
	.A0 (bus_request) );
   OAI21XL i_13 ( .Y (n_33),
	.B0 (n_49),
	.A1 (n_34),
	.A0 (n_31) );
   NAND2X1 i_2 ( .Y (n_34),
	.B (tdsp_state[1]),
	.A (tdsp_state[2]) );
   NOR2BX1 i_1 ( .Y (n_35),
	.B (tdsp_state[2]),
	.AN (tdsp_state[1]) );
   NOR2BX1 i_08999 ( .Y (n_36),
	.B (bus_grant),
	.AN (bus_request) );
   NOR2X1 i_9 ( .Y (n_37),
	.B (tdsp_state[0]),
	.A (n_36) );
   NOR2X1 i_4 ( .Y (n_40),
	.B (tdsp_state[0]),
	.A (tdsp_state[1]) );
   NAND4BXL i_17 ( .Y (n_45),
	.D (n_42),
	.C (n_102),
	.B (n_117),
	.AN (n_57) );
   AOI22X1 i_24 ( .Y (n_47),
	.B1 (n_2818),
	.B0 (tdsp_state[2]),
	.A1 (n_36),
	.A0 (n_35) );
   NOR2X1 i_35 ( .Y (n_48),
	.B (tdsp_state[2]),
	.A (n_36) );
   SDFFRHQX1 tdsp_state_reg_0 ( .SI (BG_scan_in),
	.SE (scan_en),
	.RN (n_2820),
	.Q (tdsp_state[0]),
	.D (n_33),
	.CK (clk) );
   SDFFRHQX1 tdsp_state_reg_1 ( .SI (tdsp_state[0]),
	.SE (scan_en),
	.RN (n_2820),
	.Q (tdsp_state[1]),
	.D (n_28),
	.CK (clk) );
   SDFFRHQX1 tdsp_state_reg_2 ( .SI (tdsp_state[1]),
	.SE (scan_en),
	.RN (n_2820),
	.Q (tdsp_state[2]),
	.D (n_27),
	.CK (clk) );
   SDFFHQX1 samp_bio_reg ( .SI (tdsp_state[2]),
	.SE (scan_en),
	.Q (samp_bio),
	.D (bio),
	.CK (clk) );
   SDFFHQX1 samp_int_reg ( .SI (samp_bio),
	.SE (scan_en),
	.Q (samp_int),
	.D (int),
	.CK (clk) );
   SDFFRHQX1 phi_5_reg ( .SI (samp_int),
	.SE (scan_en),
	.RN (n_2820),
	.Q (phi_5),
	.D (n_2782),
	.CK (clk) );
   OAI21XL i_598 ( .Y (n_2782),
	.B0 (n_2784),
	.A1 (n_2822),
	.A0 (n_24) );
   NAND3X1 i_599 ( .Y (n_2784),
	.C (n_24),
	.B (n_40),
	.A (tdsp_state[2]) );
   AOI21X1 i_37 ( .Y (n_49),
	.B0 (n_40),
	.A1 (n_2818),
	.A0 (n_48) );
   SDFFRHQX1 phi_4_reg ( .SI (phi_5),
	.SE (scan_en),
	.RN (n_2820),
	.Q (phi_4),
	.D (n_2788),
	.CK (clk) );
   OAI21XL i_605 ( .Y (n_2788),
	.B0 (n_2790),
	.A1 (n_2821),
	.A0 (n_24) );
   NAND3X1 i_606 ( .Y (n_2790),
	.C (n_24),
	.B (n_35),
	.A (tdsp_state[0]) );
   NOR3X1 i_20 ( .Y (n_57),
	.C (tdsp_state[0]),
	.B (tdsp_state[2]),
	.A (tdsp_state[1]) );
   SDFFRHQX1 phi_3_reg ( .SI (phi_4),
	.SE (scan_en),
	.RN (n_2820),
	.Q (phi_3),
	.D (n_2794),
	.CK (clk) );
   OAI21XL i_612 ( .Y (n_2794),
	.B0 (n_2797),
	.A1 (n_2819),
	.A0 (n_22) );
   NAND2X1 i_614 ( .Y (n_2797),
	.B (n_2819),
	.A (phi_3) );
   OR3XL i_23 ( .Y (n_72),
	.C (n_2818),
	.B (tdsp_state[1]),
	.A (tdsp_state[2]) );
   SDFFRHQX1 phi_2_reg ( .SI (phi_3),
	.SE (scan_en),
	.RN (n_2820),
	.Q (phi_2),
	.D (n_2800),
	.CK (clk) );
   OAI21XL i_619 ( .Y (n_2800),
	.B0 (n_2803),
	.A1 (n_2819),
	.A0 (n_72) );
   NAND2X1 i_621 ( .Y (n_2803),
	.B (n_2819),
	.A (phi_2) );
   NAND2X1 i_31 ( .Y (n_102),
	.B (tdsp_state[0]),
	.A (n_35) );
   SDFFRHQX1 phi_1_reg ( .SI (phi_2),
	.SE (scan_en),
	.RN (n_2820),
	.Q (phi_1),
	.D (n_2806),
	.CK (clk) );
   MX2X1 i_626 ( .Y (n_2806),
	.S0 (n_2819),
	.B (phi_1),
	.A (n_57) );
   NAND2X1 i_34 ( .Y (n_117),
	.B (n_40),
	.A (tdsp_state[2]) );
   SDFFRHQX1 phi_6_reg ( .SI (phi_1),
	.SE (scan_en),
	.RN (n_2820),
	.Q (BG_scan_out),
	.D (n_2812),
	.CK (clk) );
   OAI21XL i_633 ( .Y (n_2812),
	.B0 (n_2815),
	.A1 (n_2819),
	.A0 (n_42) );
   NAND2X1 i_635 ( .Y (n_2815),
	.B (n_2819),
	.A (phi_6) );
   NAND3BX1 i_36 ( .Y (n_42),
	.C (tdsp_state[0]),
	.B (tdsp_state[2]),
	.AN (tdsp_state[1]) );
   INVX1 i_682 ( .Y (n_2818),
	.A (tdsp_state[0]) );
   INVX1 i_683 ( .Y (n_2819),
	.A (n_24) );
   INVX1 i_684 ( .Y (n_2820),
	.A (reset) );
   INVX1 i_685 ( .Y (n_2821),
	.A (phi_4) );
   INVX1 i_686 ( .Y (n_2822),
	.A (phi_5) );
endmodule

module tdsp_core (
	clk,
	reset,
	as,
	read,
	write,
	address,
	t_data_in,
	t_data_out,
	p_read,
	p_address,
	rom_data_in,
	bus_grant,
	bus_request,
	port_as,
	port_address,
	port_pad_data_in,
	port_pad_data_out,
	bio,
	int,
	scan_en,
	BG_scan_in,
	BG_scan_out );
   input clk;
   input reset;
   output as;
   output read;
   output write;
   output [7:0] address;
   input [15:0] t_data_in;
   output [15:0] t_data_out;
   output p_read;
   output [8:0] p_address;
   input [15:0] rom_data_in;
   input bus_grant;
   output bus_request;
   output port_as;
   output [2:0] port_address;
   input [15:0] port_pad_data_in;
   output [15:0] port_pad_data_out;
   input bio;
   input int;
   input scan_en;
   input BG_scan_in;
   output BG_scan_out;

   // Internal wires
   wire [15:0] data_out;
   wire [15:0] data_in;
   wire [15:0] ir;
   wire [15:0] port_data_in;
   wire [2:0] port_addrs_in;
   wire [8:0] p_addrs_in;
   wire [2:0] sel_op_b;
   wire [2:0] sel_op_a;
   wire [15:0] top;
   wire [31:0] p;
   wire [15:0] ar1;
   wire [15:0] ar0;
   wire [15:0] port_data_out;
   wire [15:0] p_data_out;
   wire [7:0] addrs_in;
   wire [15:0] decode;
   wire [15:0] ar;
   wire [15:0] mdr;
   wire [31:0] mpy_result;
   wire [32:0] alu_result;
   wire [3:0] alu_cmd;
   wire [31:0] opb;
   wire [31:0] opa;
   wire samp_bio;
   wire phi_1;
   wire phi_3;
   wire phi_4;
   wire phi_5;
   wire phi_6;
   wire n_7866;
   wire read_prog;
   wire go_prog;
   wire n_7867;
   wire read_port;
   wire go_port;
   wire n_7868;
   wire ovm;
   wire UNCONNECTED_000;
   wire \acc[31] ;
   wire \acc[30] ;
   wire \acc[29] ;
   wire \acc[28] ;
   wire \acc[27] ;
   wire \acc[26] ;
   wire \acc[25] ;
   wire \acc[24] ;
   wire \acc[23] ;
   wire \acc[22] ;
   wire \acc[21] ;
   wire \acc[20] ;
   wire \acc[19] ;
   wire \acc[18] ;
   wire \acc[17] ;
   wire \acc[16] ;
   wire \acc[15] ;
   wire \acc[14] ;
   wire \acc[13] ;
   wire \acc[12] ;
   wire \acc[11] ;
   wire \acc[10] ;
   wire \acc[9] ;
   wire \acc[8] ;
   wire \acc[7] ;
   wire \acc[6] ;
   wire \acc[5] ;
   wire \acc[4] ;
   wire \acc[3] ;
   wire \acc[2] ;
   wire \acc[1] ;
   wire \acc[0] ;
   wire gez;
   wire gz;
   wire nz;
   wire lz;
   wire lez;
   wire arnz;
   wire bioz;
   wire skip_one;
   wire pc_acc;
   wire dmov_inc;
   wire dp;
   wire arp;
   wire UNCONNECTED_001;
   wire UNCONNECTED_002;
   wire UNCONNECTED_003;
   wire UNCONNECTED_004;
   wire UNCONNECTED_005;
   wire UNCONNECTED_006;
   wire UNCONNECTED_007;
   wire \pc[8] ;
   wire \pc[7] ;
   wire \pc[6] ;
   wire \pc[5] ;
   wire \pc[4] ;
   wire \pc[3] ;
   wire \pc[2] ;
   wire \pc[1] ;
   wire \pc[0] ;
   wire UNCONNECTED_008;
   wire enc_read_prog;
   wire enc_go_prog;
   wire enc_read_data;
   wire enc_go_data;
   wire enc_read_port;
   wire enc_go_port;
   wire n_7869;
   wire dec_read_prog;
   wire dec_go_prog;
   wire dec_read_data;
   wire dec_go_data;
   wire dec_read_port;
   wire dec_go_port;
   wire n_7870;
   wire go_data;
   wire read_data;
   wire UNCONNECTED_009;
   wire UNCONNECTED_010;
   wire UNCONNECTED_011;
   wire UNCONNECTED_012;
   wire UNCONNECTED_013;
   wire UNCONNECTED_014;
   wire UNCONNECTED_015;
   wire UNCONNECTED_016;

   tdsp_core_mach TDSP_CORE_MACH_INST ( .samp_bio (samp_bio),
	.phi_1 (phi_1),
	.phi_3 (phi_3),
	.phi_4 (phi_4),
	.phi_5 (phi_5),
	.phi_6 (phi_6),
	.reset (reset),
	.clk (clk),
	.bus_request (bus_request),
	.bus_grant (bus_grant),
	.bio (bio),
	.int (int),
	.scan_en (scan_en),
	.BG_scan_in (BG_scan_in),
	.BG_scan_out (n_7866) );
   prog_bus_mach PROG_BUS_MACH_INST ( .clk (clk),
	.reset (reset),
	.read (p_read),
	.address ({ p_address[8],
		p_address[7],
		p_address[6],
		p_address[5],
		p_address[4],
		p_address[3],
		p_address[2],
		p_address[1],
		p_address[0] }),
	.data_out ({ p_data_out[15],
		p_data_out[14],
		p_data_out[13],
		p_data_out[12],
		p_data_out[11],
		p_data_out[10],
		p_data_out[9],
		p_data_out[8],
		p_data_out[7],
		p_data_out[6],
		p_data_out[5],
		p_data_out[4],
		p_data_out[3],
		p_data_out[2],
		p_data_out[1],
		p_data_out[0] }),
	.pad_data_in ({ rom_data_in[15],
		rom_data_in[14],
		rom_data_in[13],
		rom_data_in[12],
		rom_data_in[11],
		rom_data_in[10],
		rom_data_in[9],
		rom_data_in[8],
		rom_data_in[7],
		rom_data_in[6],
		rom_data_in[5],
		rom_data_in[4],
		rom_data_in[3],
		rom_data_in[2],
		rom_data_in[1],
		rom_data_in[0] }),
	.addrs_in ({ p_addrs_in[8],
		p_addrs_in[7],
		p_addrs_in[6],
		p_addrs_in[5],
		p_addrs_in[4],
		p_addrs_in[3],
		p_addrs_in[2],
		p_addrs_in[1],
		p_addrs_in[0] }),
	.read_cycle (read_prog),
	.go (go_prog),
	.scan_en (scan_en),
	.BG_scan_in (n_7866),
	.BG_scan_out (n_7867) );
   port_bus_mach PORT_BUS_MACH_INST ( .clk (clk),
	.reset (reset),
	.address ({ port_address[2],
		port_address[1],
		port_address[0] }),
	.data_in ({ port_data_in[15],
		port_data_in[14],
		port_data_in[13],
		port_data_in[12],
		port_data_in[11],
		port_data_in[10],
		port_data_in[9],
		port_data_in[8],
		port_data_in[7],
		port_data_in[6],
		port_data_in[5],
		port_data_in[4],
		port_data_in[3],
		port_data_in[2],
		port_data_in[1],
		port_data_in[0] }),
	.data_out ({ port_data_out[15],
		port_data_out[14],
		port_data_out[13],
		port_data_out[12],
		port_data_out[11],
		port_data_out[10],
		port_data_out[9],
		port_data_out[8],
		port_data_out[7],
		port_data_out[6],
		port_data_out[5],
		port_data_out[4],
		port_data_out[3],
		port_data_out[2],
		port_data_out[1],
		port_data_out[0] }),
	.pad_data_in ({ port_pad_data_in[15],
		port_pad_data_in[14],
		port_pad_data_in[13],
		port_pad_data_in[12],
		port_pad_data_in[11],
		port_pad_data_in[10],
		port_pad_data_in[9],
		port_pad_data_in[8],
		port_pad_data_in[7],
		port_pad_data_in[6],
		port_pad_data_in[5],
		port_pad_data_in[4],
		port_pad_data_in[3],
		port_pad_data_in[2],
		port_pad_data_in[1],
		port_pad_data_in[0] }),
	.pad_data_out ({ port_pad_data_out[15],
		port_pad_data_out[14],
		port_pad_data_out[13],
		port_pad_data_out[12],
		port_pad_data_out[11],
		port_pad_data_out[10],
		port_pad_data_out[9],
		port_pad_data_out[8],
		port_pad_data_out[7],
		port_pad_data_out[6],
		port_pad_data_out[5],
		port_pad_data_out[4],
		port_pad_data_out[3],
		port_pad_data_out[2],
		port_pad_data_out[1],
		port_pad_data_out[0] }),
	.addrs_in ({ port_addrs_in[2],
		port_addrs_in[1],
		port_addrs_in[0] }),
	.read_cycle (read_port),
	.go (go_port),
	.as (port_as),
	.scan_en (scan_en),
	.BG_scan_in (n_7867),
	.BG_scan_out (n_7868) );
   alu_32 ALU_32_INST ( .ovm (ovm),
	.op_a ({ opa[31],
		opa[30],
		opa[29],
		opa[28],
		opa[27],
		opa[26],
		opa[25],
		opa[24],
		opa[23],
		opa[22],
		opa[21],
		opa[20],
		opa[19],
		opa[18],
		opa[17],
		opa[16],
		opa[15],
		opa[14],
		opa[13],
		opa[12],
		opa[11],
		opa[10],
		opa[9],
		opa[8],
		opa[7],
		opa[6],
		opa[5],
		opa[4],
		opa[3],
		opa[2],
		opa[1],
		opa[0] }),
	.op_b ({ opb[31],
		opb[30],
		opb[29],
		opb[28],
		opb[27],
		opb[26],
		opb[25],
		opb[24],
		opb[23],
		opb[22],
		opb[21],
		opb[20],
		opb[19],
		opb[18],
		opb[17],
		opb[16],
		opb[15],
		opb[14],
		opb[13],
		opb[12],
		opb[11],
		opb[10],
		opb[9],
		opb[8],
		opb[7],
		opb[6],
		opb[5],
		opb[4],
		opb[3],
		opb[2],
		opb[1],
		opb[0] }),
	.result ({ alu_result[32],
		alu_result[31],
		alu_result[30],
		alu_result[29],
		alu_result[28],
		alu_result[27],
		alu_result[26],
		alu_result[25],
		alu_result[24],
		alu_result[23],
		alu_result[22],
		alu_result[21],
		alu_result[20],
		alu_result[19],
		alu_result[18],
		alu_result[17],
		alu_result[16],
		alu_result[15],
		alu_result[14],
		alu_result[13],
		alu_result[12],
		alu_result[11],
		alu_result[10],
		alu_result[9],
		alu_result[8],
		alu_result[7],
		alu_result[6],
		alu_result[5],
		alu_result[4],
		alu_result[3],
		alu_result[2],
		alu_result[1],
		alu_result[0] }),
	.cmd ({ alu_cmd[3],
		alu_cmd[2],
		alu_cmd[1],
		alu_cmd[0] }) );
   mult_32 MPY_32_INST ( .op_a ({ opa[15],
		opa[14],
		opa[13],
		opa[12],
		opa[11],
		opa[10],
		opa[9],
		opa[8],
		opa[7],
		opa[6],
		opa[5],
		opa[4],
		opa[3],
		opa[2],
		opa[1],
		opa[0] }),
	.op_b ({ opb[15],
		opb[14],
		opb[13],
		opb[12],
		opb[11],
		opb[10],
		opb[9],
		opb[8],
		opb[7],
		opb[6],
		opb[5],
		opb[4],
		opb[3],
		opb[2],
		opb[1],
		opb[0] }),
	.result ({ mpy_result[31],
		mpy_result[30],
		mpy_result[29],
		mpy_result[28],
		mpy_result[27],
		mpy_result[26],
		mpy_result[25],
		mpy_result[24],
		mpy_result[23],
		mpy_result[22],
		mpy_result[21],
		mpy_result[20],
		mpy_result[19],
		mpy_result[18],
		mpy_result[17],
		mpy_result[16],
		mpy_result[15],
		mpy_result[14],
		mpy_result[13],
		mpy_result[12],
		mpy_result[11],
		mpy_result[10],
		mpy_result[9],
		mpy_result[8],
		mpy_result[7],
		mpy_result[6],
		mpy_result[5],
		mpy_result[4],
		mpy_result[3],
		mpy_result[2],
		mpy_result[1],
		mpy_result[0] }) );
   accum_stat ACCUM_STAT_INST ( .accum ({ UNCONNECTED_000,
		\acc[31] ,
		\acc[30] ,
		\acc[29] ,
		\acc[28] ,
		\acc[27] ,
		\acc[26] ,
		\acc[25] ,
		\acc[24] ,
		\acc[23] ,
		\acc[22] ,
		\acc[21] ,
		\acc[20] ,
		\acc[19] ,
		\acc[18] ,
		\acc[17] ,
		\acc[16] ,
		\acc[15] ,
		\acc[14] ,
		\acc[13] ,
		\acc[12] ,
		\acc[11] ,
		\acc[10] ,
		\acc[9] ,
		\acc[8] ,
		\acc[7] ,
		\acc[6] ,
		\acc[5] ,
		\acc[4] ,
		\acc[3] ,
		\acc[2] ,
		\acc[1] ,
		\acc[0]  }),
	.ar ({ ar[15],
		ar[14],
		ar[13],
		ar[12],
		ar[11],
		ar[10],
		ar[9],
		ar[8],
		ar[7],
		ar[6],
		ar[5],
		ar[4],
		ar[3],
		ar[2],
		ar[1],
		ar[0] }),
	.bio (samp_bio),
	.gez (gez),
	.gz (gz),
	.nz (nz),
	.lz (lz),
	.lez (lez),
	.arnz (arnz),
	.bioz (bioz) );
   execute_i EXECUTE_INST ( .clk (clk),
	.reset (reset),
	.phi_1 (phi_1),
	.phi_3 (phi_3),
	.phi_4 (phi_4),
	.phi_5 (phi_5),
	.phi_6 (phi_6),
	.gez (gez),
	.gz (gz),
	.nz (nz),
	.lz (lz),
	.lez (lez),
	.arnz (arnz),
	.bioz (bioz),
	.alu_result ({ alu_result[32],
		alu_result[31],
		alu_result[30],
		alu_result[29],
		alu_result[28],
		alu_result[27],
		alu_result[26],
		alu_result[25],
		alu_result[24],
		alu_result[23],
		alu_result[22],
		alu_result[21],
		alu_result[20],
		alu_result[19],
		alu_result[18],
		alu_result[17],
		alu_result[16],
		alu_result[15],
		alu_result[14],
		alu_result[13],
		alu_result[12],
		alu_result[11],
		alu_result[10],
		alu_result[9],
		alu_result[8],
		alu_result[7],
		alu_result[6],
		alu_result[5],
		alu_result[4],
		alu_result[3],
		alu_result[2],
		alu_result[1],
		alu_result[0] }),
	.mpy_result ({ mpy_result[31],
		mpy_result[30],
		mpy_result[29],
		mpy_result[28],
		mpy_result[27],
		mpy_result[26],
		mpy_result[25],
		mpy_result[24],
		mpy_result[23],
		mpy_result[22],
		mpy_result[21],
		mpy_result[20],
		mpy_result[19],
		mpy_result[18],
		mpy_result[17],
		mpy_result[16],
		mpy_result[15],
		mpy_result[14],
		mpy_result[13],
		mpy_result[12],
		mpy_result[11],
		mpy_result[10],
		mpy_result[9],
		mpy_result[8],
		mpy_result[7],
		mpy_result[6],
		mpy_result[5],
		mpy_result[4],
		mpy_result[3],
		mpy_result[2],
		mpy_result[1],
		mpy_result[0] }),
	.mdr ({ mdr[15],
		mdr[14],
		mdr[13],
		mdr[12],
		mdr[11],
		mdr[10],
		mdr[9],
		mdr[8],
		mdr[7],
		mdr[6],
		mdr[5],
		mdr[4],
		mdr[3],
		mdr[2],
		mdr[1],
		mdr[0] }),
	.ir ({ ir[15],
		ir[14],
		ir[13],
		ir[12],
		ir[11],
		ir[10],
		ir[9],
		ir[8],
		ir[7],
		ir[6],
		ir[5],
		ir[4],
		ir[3],
		ir[2],
		ir[1],
		ir[0] }),
	.decode ({ decode[15],
		decode[14],
		decode[13],
		decode[12],
		decode[11],
		decode[10],
		decode[9],
		decode[8],
		decode[7],
		decode[6],
		decode[5],
		decode[4],
		decode[3],
		decode[2],
		decode[1],
		decode[0] }),
	.ar ({ ar[15],
		ar[14],
		ar[13],
		ar[12],
		ar[11],
		ar[10],
		ar[9],
		ar[8],
		ar[7],
		ar[6],
		ar[5],
		ar[4],
		ar[3],
		ar[2],
		ar[1],
		ar[0] }),
	.skip_one (skip_one),
	.pc_acc (pc_acc),
	.dmov_inc (dmov_inc),
	.dp (dp),
	.arp (arp),
	.ar0 ({ ar0[15],
		ar0[14],
		ar0[13],
		ar0[12],
		ar0[11],
		ar0[10],
		ar0[9],
		ar0[8],
		ar0[7],
		ar0[6],
		ar0[5],
		ar0[4],
		ar0[3],
		ar0[2],
		ar0[1],
		ar0[0] }),
	.ar1 ({ ar1[15],
		ar1[14],
		ar1[13],
		ar1[12],
		ar1[11],
		ar1[10],
		ar1[9],
		ar1[8],
		ar1[7],
		ar1[6],
		ar1[5],
		ar1[4],
		ar1[3],
		ar1[2],
		ar1[1],
		ar1[0] }),
	.pc ({ UNCONNECTED_001,
		UNCONNECTED_002,
		UNCONNECTED_003,
		UNCONNECTED_004,
		UNCONNECTED_005,
		UNCONNECTED_006,
		UNCONNECTED_007,
		\pc[8] ,
		\pc[7] ,
		\pc[6] ,
		\pc[5] ,
		\pc[4] ,
		\pc[3] ,
		\pc[2] ,
		\pc[1] ,
		\pc[0]  }),
	.acc ({ UNCONNECTED_008,
		\acc[31] ,
		\acc[30] ,
		\acc[29] ,
		\acc[28] ,
		\acc[27] ,
		\acc[26] ,
		\acc[25] ,
		\acc[24] ,
		\acc[23] ,
		\acc[22] ,
		\acc[21] ,
		\acc[20] ,
		\acc[19] ,
		\acc[18] ,
		\acc[17] ,
		\acc[16] ,
		\acc[15] ,
		\acc[14] ,
		\acc[13] ,
		\acc[12] ,
		\acc[11] ,
		\acc[10] ,
		\acc[9] ,
		\acc[8] ,
		\acc[7] ,
		\acc[6] ,
		\acc[5] ,
		\acc[4] ,
		\acc[3] ,
		\acc[2] ,
		\acc[1] ,
		\acc[0]  }),
	.p ({ p[31],
		p[30],
		p[29],
		p[28],
		p[27],
		p[26],
		p[25],
		p[24],
		p[23],
		p[22],
		p[21],
		p[20],
		p[19],
		p[18],
		p[17],
		p[16],
		p[15],
		p[14],
		p[13],
		p[12],
		p[11],
		p[10],
		p[9],
		p[8],
		p[7],
		p[6],
		p[5],
		p[4],
		p[3],
		p[2],
		p[1],
		p[0] }),
	.top ({ top[15],
		top[14],
		top[13],
		top[12],
		top[11],
		top[10],
		top[9],
		top[8],
		top[7],
		top[6],
		top[5],
		top[4],
		top[3],
		top[2],
		top[1],
		top[0] }),
	.alu_cmd ({ alu_cmd[3],
		alu_cmd[2],
		alu_cmd[1],
		alu_cmd[0] }),
	.sel_op_a ({ sel_op_a[2],
		sel_op_a[1],
		sel_op_a[0] }),
	.sel_op_b ({ sel_op_b[2],
		sel_op_b[1],
		sel_op_b[0] }),
	.read_prog (enc_read_prog),
	.go_prog (enc_go_prog),
	.read_data (enc_read_data),
	.go_data (enc_go_data),
	.read_port (enc_read_port),
	.go_port (enc_go_port),
	.ovm (ovm),
	.scan_en (scan_en),
	.BG_scan_in (n_7868),
	.BG_scan_out (n_7869) );
   decode_i DECODE_INST ( .clk (clk),
	.reset (reset),
	.phi_3 (phi_3),
	.phi_6 (phi_6),
	.decode ({ decode[15],
		decode[14],
		decode[13],
		decode[12],
		decode[11],
		decode[10],
		decode[9],
		decode[8],
		decode[7],
		decode[6],
		decode[5],
		decode[4],
		decode[3],
		decode[2],
		decode[1],
		decode[0] }),
	.p_data_out ({ p_data_out[15],
		p_data_out[14],
		p_data_out[13],
		p_data_out[12],
		p_data_out[11],
		p_data_out[10],
		p_data_out[9],
		p_data_out[8],
		p_data_out[7],
		p_data_out[6],
		p_data_out[5],
		p_data_out[4],
		p_data_out[3],
		p_data_out[2],
		p_data_out[1],
		p_data_out[0] }),
	.ir ({ ir[15],
		ir[14],
		ir[13],
		ir[12],
		ir[11],
		ir[10],
		ir[9],
		ir[8],
		ir[7],
		ir[6],
		ir[5],
		ir[4],
		ir[3],
		ir[2],
		ir[1],
		ir[0] }),
	.skip_one (skip_one),
	.read_prog (dec_read_prog),
	.go_prog (dec_go_prog),
	.read_data (dec_read_data),
	.go_data (dec_go_data),
	.read_port (dec_read_port),
	.go_port (dec_go_port),
	.scan_en (scan_en),
	.BG_scan_in (n_7869),
	.BG_scan_out (n_7870) );
   tdsp_core_glue TDSP_CORE_GLUE_INST ( .addrs_in ({ addrs_in[7],
		addrs_in[6],
		addrs_in[5],
		addrs_in[4],
		addrs_in[3],
		addrs_in[2],
		addrs_in[1],
		addrs_in[0] }),
	.data_in ({ data_in[15],
		data_in[14],
		data_in[13],
		data_in[12],
		data_in[11],
		data_in[10],
		data_in[9],
		data_in[8],
		data_in[7],
		data_in[6],
		data_in[5],
		data_in[4],
		data_in[3],
		data_in[2],
		data_in[1],
		data_in[0] }),
	.p_addrs_in ({ p_addrs_in[8],
		p_addrs_in[7],
		p_addrs_in[6],
		p_addrs_in[5],
		p_addrs_in[4],
		p_addrs_in[3],
		p_addrs_in[2],
		p_addrs_in[1],
		p_addrs_in[0] }),
	.port_addrs_in ({ port_addrs_in[2],
		port_addrs_in[1],
		port_addrs_in[0] }),
	.port_data_in ({ port_data_in[15],
		port_data_in[14],
		port_data_in[13],
		port_data_in[12],
		port_data_in[11],
		port_data_in[10],
		port_data_in[9],
		port_data_in[8],
		port_data_in[7],
		port_data_in[6],
		port_data_in[5],
		port_data_in[4],
		port_data_in[3],
		port_data_in[2],
		port_data_in[1],
		port_data_in[0] }),
	.ar ({ ar[15],
		ar[14],
		ar[13],
		ar[12],
		ar[11],
		ar[10],
		ar[9],
		ar[8],
		ar[7],
		ar[6],
		ar[5],
		ar[4],
		ar[3],
		ar[2],
		ar[1],
		ar[0] }),
	.go_prog (go_prog),
	.read_prog (read_prog),
	.go_data (go_data),
	.read_data (read_data),
	.go_port (go_port),
	.read_port (read_port),
	.pc_acc (pc_acc),
	.arp (arp),
	.ar1 ({ ar1[15],
		ar1[14],
		ar1[13],
		ar1[12],
		ar1[11],
		ar1[10],
		ar1[9],
		ar1[8],
		ar1[7],
		ar1[6],
		ar1[5],
		ar1[4],
		ar1[3],
		ar1[2],
		ar1[1],
		ar1[0] }),
	.ar0 ({ ar0[15],
		ar0[14],
		ar0[13],
		ar0[12],
		ar0[11],
		ar0[10],
		ar0[9],
		ar0[8],
		ar0[7],
		ar0[6],
		ar0[5],
		ar0[4],
		ar0[3],
		ar0[2],
		ar0[1],
		ar0[0] }),
	.dp (dp),
	.ir ({ ir[15],
		ir[14],
		ir[13],
		ir[12],
		ir[11],
		ir[10],
		ir[9],
		ir[8],
		ir[7],
		ir[6],
		ir[5],
		ir[4],
		ir[3],
		ir[2],
		ir[1],
		ir[0] }),
	.opa ({ opa[31],
		opa[30],
		opa[29],
		opa[28],
		opa[27],
		opa[26],
		opa[25],
		opa[24],
		opa[23],
		opa[22],
		opa[21],
		opa[20],
		opa[19],
		opa[18],
		opa[17],
		opa[16],
		opa[15],
		opa[14],
		opa[13],
		opa[12],
		opa[11],
		opa[10],
		opa[9],
		opa[8],
		opa[7],
		opa[6],
		opa[5],
		opa[4],
		opa[3],
		opa[2],
		opa[1],
		opa[0] }),
	.opb ({ opb[31],
		opb[30],
		opb[29],
		opb[28],
		opb[27],
		opb[26],
		opb[25],
		opb[24],
		opb[23],
		opb[22],
		opb[21],
		opb[20],
		opb[19],
		opb[18],
		opb[17],
		opb[16],
		opb[15],
		opb[14],
		opb[13],
		opb[12],
		opb[11],
		opb[10],
		opb[9],
		opb[8],
		opb[7],
		opb[6],
		opb[5],
		opb[4],
		opb[3],
		opb[2],
		opb[1],
		opb[0] }),
	.mdr ({ mdr[15],
		mdr[14],
		mdr[13],
		mdr[12],
		mdr[11],
		mdr[10],
		mdr[9],
		mdr[8],
		mdr[7],
		mdr[6],
		mdr[5],
		mdr[4],
		mdr[3],
		mdr[2],
		mdr[1],
		mdr[0] }),
	.acc ({ UNCONNECTED_009,
		\acc[31] ,
		\acc[30] ,
		\acc[29] ,
		\acc[28] ,
		\acc[27] ,
		\acc[26] ,
		\acc[25] ,
		\acc[24] ,
		\acc[23] ,
		\acc[22] ,
		\acc[21] ,
		\acc[20] ,
		\acc[19] ,
		\acc[18] ,
		\acc[17] ,
		\acc[16] ,
		\acc[15] ,
		\acc[14] ,
		\acc[13] ,
		\acc[12] ,
		\acc[11] ,
		\acc[10] ,
		\acc[9] ,
		\acc[8] ,
		\acc[7] ,
		\acc[6] ,
		\acc[5] ,
		\acc[4] ,
		\acc[3] ,
		\acc[2] ,
		\acc[1] ,
		\acc[0]  }),
	.pc ({ UNCONNECTED_010,
		UNCONNECTED_011,
		UNCONNECTED_012,
		UNCONNECTED_013,
		UNCONNECTED_014,
		UNCONNECTED_015,
		UNCONNECTED_016,
		\pc[8] ,
		\pc[7] ,
		\pc[6] ,
		\pc[5] ,
		\pc[4] ,
		\pc[3] ,
		\pc[2] ,
		\pc[1] ,
		\pc[0]  }),
	.data_out ({ data_out[15],
		data_out[14],
		data_out[13],
		data_out[12],
		data_out[11],
		data_out[10],
		data_out[9],
		data_out[8],
		data_out[7],
		data_out[6],
		data_out[5],
		data_out[4],
		data_out[3],
		data_out[2],
		data_out[1],
		data_out[0] }),
	.p_data_out ({ p_data_out[15],
		p_data_out[14],
		p_data_out[13],
		p_data_out[12],
		p_data_out[11],
		p_data_out[10],
		p_data_out[9],
		p_data_out[8],
		p_data_out[7],
		p_data_out[6],
		p_data_out[5],
		p_data_out[4],
		p_data_out[3],
		p_data_out[2],
		p_data_out[1],
		p_data_out[0] }),
	.port_data_out ({ port_data_out[15],
		port_data_out[14],
		port_data_out[13],
		port_data_out[12],
		port_data_out[11],
		port_data_out[10],
		port_data_out[9],
		port_data_out[8],
		port_data_out[7],
		port_data_out[6],
		port_data_out[5],
		port_data_out[4],
		port_data_out[3],
		port_data_out[2],
		port_data_out[1],
		port_data_out[0] }),
	.top ({ top[15],
		top[14],
		top[13],
		top[12],
		top[11],
		top[10],
		top[9],
		top[8],
		top[7],
		top[6],
		top[5],
		top[4],
		top[3],
		top[2],
		top[1],
		top[0] }),
	.p ({ p[31],
		p[30],
		p[29],
		p[28],
		p[27],
		p[26],
		p[25],
		p[24],
		p[23],
		p[22],
		p[21],
		p[20],
		p[19],
		p[18],
		p[17],
		p[16],
		p[15],
		p[14],
		p[13],
		p[12],
		p[11],
		p[10],
		p[9],
		p[8],
		p[7],
		p[6],
		p[5],
		p[4],
		p[3],
		p[2],
		p[1],
		p[0] }),
	.sel_op_a ({ sel_op_a[2],
		sel_op_a[1],
		sel_op_a[0] }),
	.sel_op_b ({ sel_op_b[2],
		sel_op_b[1],
		sel_op_b[0] }),
	.dec_go_prog (dec_go_prog),
	.enc_go_prog (enc_go_prog),
	.dec_read_prog (dec_read_prog),
	.enc_read_prog (enc_read_prog),
	.dec_go_data (dec_go_data),
	.enc_go_data (enc_go_data),
	.dec_read_data (dec_read_data),
	.enc_read_data (enc_read_data),
	.dec_go_port (dec_go_port),
	.enc_go_port (enc_go_port),
	.dec_read_port (dec_read_port),
	.enc_read_port (enc_read_port),
	.dmov_inc (dmov_inc) );
   data_bus_mach DATA_BUS_MACH_INST ( .clk (clk),
	.reset (reset),
	.read (read),
	.write (write),
	.address ({ address[7],
		address[6],
		address[5],
		address[4],
		address[3],
		address[2],
		address[1],
		address[0] }),
	.data_in ({ data_in[15],
		data_in[14],
		data_in[13],
		data_in[12],
		data_in[11],
		data_in[10],
		data_in[9],
		data_in[8],
		data_in[7],
		data_in[6],
		data_in[5],
		data_in[4],
		data_in[3],
		data_in[2],
		data_in[1],
		data_in[0] }),
	.data_out ({ data_out[15],
		data_out[14],
		data_out[13],
		data_out[12],
		data_out[11],
		data_out[10],
		data_out[9],
		data_out[8],
		data_out[7],
		data_out[6],
		data_out[5],
		data_out[4],
		data_out[3],
		data_out[2],
		data_out[1],
		data_out[0] }),
	.pad_data_in ({ t_data_in[15],
		t_data_in[14],
		t_data_in[13],
		t_data_in[12],
		t_data_in[11],
		t_data_in[10],
		t_data_in[9],
		t_data_in[8],
		t_data_in[7],
		t_data_in[6],
		t_data_in[5],
		t_data_in[4],
		t_data_in[3],
		t_data_in[2],
		t_data_in[1],
		t_data_in[0] }),
	.pad_data_out ({ t_data_out[15],
		t_data_out[14],
		t_data_out[13],
		t_data_out[12],
		t_data_out[11],
		t_data_out[10],
		t_data_out[9],
		t_data_out[8],
		t_data_out[7],
		t_data_out[6],
		t_data_out[5],
		t_data_out[4],
		t_data_out[3],
		t_data_out[2],
		t_data_out[1],
		t_data_out[0] }),
	.addrs_in ({ addrs_in[7],
		addrs_in[6],
		addrs_in[5],
		addrs_in[4],
		addrs_in[3],
		addrs_in[2],
		addrs_in[1],
		addrs_in[0] }),
	.read_cycle (read_data),
	.go (go_data),
	.as (as),
	.bus_request (bus_request),
	.bus_grant (bus_grant),
	.scan_en (scan_en),
	.BG_scan_in (n_7870),
	.BG_scan_out (BG_scan_out) );
endmodule


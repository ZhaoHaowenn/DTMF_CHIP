// Created on Fri Jun 14 13:52:44 2002

module accum_stat(
		accum,
		ar,
		bio,
		gez,
		gz,
		nz,
		z,
		lz,
		lez,
		ov,
		arnz,
		bioz);

	input [32:0] accum;
	input [15:0] ar;
	input bio;
	output gez;
	output gz;
	output nz;
	output z;
	output lz;
	output lez;
	input ov;
	output arnz;
	output bioz;




	INVXL i_9530(
		.A(n_6309),
		.Y(lz));

	INVXL i_9529(
		.A(accum[31]),
		.Y(n_6309));

	NOR2X1 i_4403(
		.A(lz),
		.B(n_73),
		.Y(gz));

	NOR4X1 i_43(
		.A(accum[2]),
		.B(accum[3]),
		.C(accum[0]),
		.D(accum[1]),
		.Y(n_46));

	NOR4X1 i_40(
		.A(accum[6]),
		.B(accum[7]),
		.C(accum[4]),
		.D(accum[5]),
		.Y(n_49));

	NOR4X1 i_36(
		.A(accum[10]),
		.B(accum[11]),
		.C(accum[8]),
		.D(accum[9]),
		.Y(n_53));

	NOR4X1 i_33(
		.A(accum[14]),
		.B(accum[15]),
		.C(accum[12]),
		.D(accum[13]),
		.Y(n_56));

	NAND4X1 i_45(
		.A(n_56),
		.B(n_53),
		.C(n_49),
		.D(n_46),
		.Y(n_58));

	OR4X1 i_28(
		.A(accum[18]),
		.B(accum[19]),
		.C(accum[16]),
		.D(accum[17]),
		.Y(n_61));

	NOR4X1 i_25(
		.A(accum[22]),
		.B(accum[23]),
		.C(accum[20]),
		.D(accum[21]),
		.Y(n_64));

	OR4X1 i_21(
		.A(accum[26]),
		.B(accum[27]),
		.C(accum[24]),
		.D(accum[25]),
		.Y(n_68));

	OR4X1 i_22(
		.A(accum[28]),
		.B(accum[29]),
		.C(accum[30]),
		.D(n_68),
		.Y(n_71));

	NOR4BX1 i_09004(
		.AN(n_64),
		.B(n_58),
		.C(n_61),
		.D(n_71),
		.Y(n_73));

	NOR4X1 i_13(
		.A(ar[2]),
		.B(ar[3]),
		.C(ar[0]),
		.D(ar[1]),
		.Y(n_76));

	NOR4X1 i_10(
		.A(ar[6]),
		.B(ar[7]),
		.C(ar[4]),
		.D(ar[5]),
		.Y(n_79));

	NOR4X1 i_6(
		.A(ar[10]),
		.B(ar[11]),
		.C(ar[8]),
		.D(ar[9]),
		.Y(n_83));

	NOR4X1 i_3(
		.A(ar[14]),
		.B(ar[15]),
		.C(ar[12]),
		.D(ar[13]),
		.Y(n_87));

	OAI21XL i_4401(
		.A0(lz),
		.A1(n_73),
		.B0(nz),
		.Y(gez));

	NAND2BX1 i_4406(
		.AN(lz),
		.B(n_73),
		.Y(nz));

	OR2X1 i_4405(
		.A(lz),
		.B(n_73),
		.Y(lez));

	NAND4X1 i_342308(
		.A(n_87),
		.B(n_83),
		.C(n_79),
		.D(n_76),
		.Y(arnz));

	INVX1 i_3339(
		.A(bio),
		.Y(bioz));

endmodule
module alu_32(
		ovm,
		op_a,
		op_b,
		result,
		cmd);

	input ovm;
	input [31:0] op_a;
	input [31:0] op_b;
	output [32:0] result;
	input [3:0] cmd;




	CLKBUFXL i_10254(
		.A(n_6939),
		.Y(n_7387));

	BUFX3 i_10242(
		.A(n_3062),
		.Y(n_7369));

	BUFX3 i_10232(
		.A(n_1942),
		.Y(n_7356));

	CLKBUFXL i_10228(
		.A(n_907),
		.Y(n_7350));

	CLKBUFXL i_10227(
		.A(n_907),
		.Y(n_7347));

	CLKBUFXL i_10225(
		.A(n_1716),
		.Y(n_7344));

	CLKBUFXL i_10223(
		.A(n_868),
		.Y(n_7341));

	BUFX2 i_10221(
		.A(n_6906),
		.Y(n_7338));

	CLKBUFXL i_10218(
		.A(n_6909),
		.Y(n_7335));

	CLKBUFXL i_10214(
		.A(n_1716),
		.Y(n_7329));

	CLKBUFXL i_10213(
		.A(n_3062),
		.Y(n_7326));

	CLKBUFXL i_10211(
		.A(n_1738),
		.Y(n_7323));

	BUFX3 i_10208(
		.A(n_7317),
		.Y(n_7320));

	CLKBUFX2 i_10206(
		.A(cmd[1]),
		.Y(n_7317));

	CLKBUFXL i_10203(
		.A(cmd[0]),
		.Y(n_7313));

	BUFX3 i_10194(
		.A(op_a[3]),
		.Y(n_7302));

	BUFXL i_10184(
		.A(op_a[10]),
		.Y(n_7290));

	BUFXL i_10168(
		.A(op_a[14]),
		.Y(n_7270));

	CLKBUFXL i_9954(
		.A(n_1738),
		.Y(n_6939));

	CLKBUFXL i_9937(
		.A(n_3068),
		.Y(n_6911));

	CLKBUFXL i_9936(
		.A(n_1727),
		.Y(n_6909));

	CLKBUFXL i_9934(
		.A(n_2071),
		.Y(n_6906));

	CLKBUFXL i_9933(
		.A(n_868),
		.Y(n_6904));

	CLKBUFXL i_9931(
		.A(n_1942),
		.Y(n_6901));

	CLKBUFXL i_9927(
		.A(n_3060),
		.Y(n_6894));

	CLKBUFXL i_9926(
		.A(n_3060),
		.Y(n_6893));

	NOR2X1 i_1454(
		.A(n_2382),
		.B(n_911),
		.Y(n_1618));

	AOI211X1 i_361(
		.A0(n_1830),
		.A1(n_1831),
		.B0(n_1827),
		.C0(n_1616),
		.Y(n_1617));

	NOR2X1 i_1451(
		.A(n_906),
		.B(n_1880),
		.Y(n_1616));

	NOR2X1 i_1449(
		.A(n_1936),
		.B(op_a[27]),
		.Y(n_1614));

	NAND2BX1 i_1448(
		.AN(n_949),
		.B(n_3062),
		.Y(n_1613));

	NAND3X1 i_446(
		.A(n_879),
		.B(n_1611),
		.C(n_1754),
		.Y(n_1612));

	NAND3BX1 i_1445(
		.AN(n_1806),
		.B(n_1758),
		.C(n_946),
		.Y(n_1611));

	OAI21XL i_778553(
		.A0(n_1609),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[26]));

	AOI211X1 i_1351(
		.A0(n_1598),
		.A1(n_2360),
		.B0(n_7335),
		.C0(n_2378),
		.Y(n_1609));

	OAI21XL i_261(
		.A0(n_2370),
		.A1(n_1699),
		.B0(n_1596),
		.Y(n_1600));

	AOI21X1 i_262(
		.A0(op_a[26]),
		.A1(n_2372),
		.B0(n_1589),
		.Y(n_1599));

	OAI2BB1X1 i_263(
		.A0N(n_1708),
		.A1N(n_7326),
		.B0(n_1716),
		.Y(n_1598));

	NAND2X1 i_1424(
		.A(n_1699),
		.B(n_2370),
		.Y(n_1596));

	AOI211X1 i_356(
		.A0(n_2264),
		.A1(n_2300),
		.B0(n_2299),
		.C0(n_1593),
		.Y(n_1594));

	NOR4BX1 i_1419(
		.AN(n_2300),
		.B(n_1441),
		.C(n_1395),
		.D(n_1494),
		.Y(n_1593));

	NOR2X1 i_251379(
		.A(op_b[25]),
		.B(op_a[25]),
		.Y(n_1592));

	NOR2X1 i_1416(
		.A(n_2372),
		.B(op_a[26]),
		.Y(n_1589));

	OAI211X1 i_445(
		.A0(n_2295),
		.A1(n_2259),
		.B0(n_2294),
		.C0(n_1586),
		.Y(n_1587));

	NAND4BXL i_1410(
		.AN(n_2260),
		.B(n_1485),
		.C(n_925),
		.D(n_1487),
		.Y(n_1586));

	NAND2BX1 i_577104(
		.AN(op_a[25]),
		.B(op_b[25]),
		.Y(n_1585));

	OAI21XL i_788554(
		.A0(n_1582),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[25]));

	AOI211X1 i_1342(
		.A0(n_1571),
		.A1(n_2341),
		.B0(n_7335),
		.C0(n_2358),
		.Y(n_1582));

	NOR2X1 i_1384(
		.A(n_1573),
		.B(n_3095),
		.Y(n_1579));

	AOI31X1 i_252(
		.A0(n_1566),
		.A1(n_2346),
		.A2(n_2349),
		.B0(n_1568),
		.Y(n_1573));

	AOI31X1 i_253(
		.A0(n_2285),
		.A1(op_a[25]),
		.A2(n_2351),
		.B0(n_1563),
		.Y(n_1572));

	OAI21XL i_254(
		.A0(n_2344),
		.A1(n_7323),
		.B0(n_7344),
		.Y(n_1571));

	AOI21X1 i_1375(
		.A0(n_1566),
		.A1(n_2346),
		.B0(n_2349),
		.Y(n_1568));

	AOI211X1 i_355(
		.A0(n_1835),
		.A1(n_1879),
		.B0(n_1830),
		.C0(n_1565),
		.Y(n_1567));

	NAND3BX1 i_1373(
		.AN(n_1567),
		.B(n_1881),
		.C(n_1831),
		.Y(n_1566));

	NOR4BX1 i_1371(
		.AN(n_1879),
		.B(n_1395),
		.C(n_1390),
		.D(n_1467),
		.Y(n_1565));

	AOI21X1 i_1368(
		.A0(n_2351),
		.A1(n_2285),
		.B0(op_a[25]),
		.Y(n_1563));

	OAI211X1 i_444(
		.A0(n_1806),
		.A1(n_1762),
		.B0(n_1757),
		.C0(n_1559),
		.Y(n_1561));

	NAND4BXL i_1361(
		.AN(n_1806),
		.B(n_1462),
		.C(n_927),
		.D(n_1383),
		.Y(n_1559));

	OAI21XL i_798555(
		.A0(n_1557),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[24]));

	AOI211X1 i_1333(
		.A0(n_1546),
		.A1(n_2323),
		.B0(n_7335),
		.C0(n_2339),
		.Y(n_1557));

	OAI21XL i_245(
		.A0(n_2333),
		.A1(n_1647),
		.B0(n_1543),
		.Y(n_1548));

	AOI21X1 i_246(
		.A0(op_a[24]),
		.A1(n_1907),
		.B0(n_1536),
		.Y(n_1547));

	OAI2BB1X1 i_248(
		.A0N(n_1637),
		.A1N(n_7326),
		.B0(n_1716),
		.Y(n_1546));

	NOR2X1 i_241378(
		.A(op_b[24]),
		.B(op_a[24]),
		.Y(n_1544));

	NAND2X1 i_1338(
		.A(n_1647),
		.B(n_2333),
		.Y(n_1543));

	AOI211X1 i_354(
		.A0(n_2233),
		.A1(n_2265),
		.B0(n_2264),
		.C0(n_1540),
		.Y(n_1541));

	NOR4BX1 i_1332(
		.AN(n_2234),
		.B(n_1441),
		.C(n_1395),
		.D(n_1443),
		.Y(n_1540));

	NOR2X1 i_231377(
		.A(op_b[23]),
		.B(op_a[23]),
		.Y(n_1539));

	NOR2X1 i_1329(
		.A(n_1907),
		.B(op_a[24]),
		.Y(n_1536));

	OAI211X1 i_437(
		.A0(n_2228),
		.A1(n_2260),
		.B0(n_2259),
		.C0(n_1533),
		.Y(n_1534));

	NAND4BXL i_1323(
		.AN(n_2260),
		.B(n_1383),
		.C(n_1436),
		.D(n_929),
		.Y(n_1533));

	NAND2BX1 i_557102(
		.AN(op_a[23]),
		.B(op_b[23]),
		.Y(n_1532));

	OAI21XL i_808556(
		.A0(n_1529),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[23]));

	AOI211X1 i_1324(
		.A0(n_1518),
		.A1(n_2313),
		.B0(n_6909),
		.C0(n_2321),
		.Y(n_1529));

	OAI21XL i_238(
		.A0(n_2315),
		.A1(n_1617),
		.B0(n_1516),
		.Y(n_1520));

	AOI31X1 i_240(
		.A0(n_1930),
		.A1(op_a[23]),
		.A2(n_1932),
		.B0(n_1513),
		.Y(n_1519));

	OAI2BB1X1 i_241(
		.A0N(n_1612),
		.A1N(n_7326),
		.B0(n_7344),
		.Y(n_1518));

	NAND2X1 i_1300(
		.A(n_1617),
		.B(n_2315),
		.Y(n_1516));

	AOI21X1 i_1296(
		.A0(n_1932),
		.A1(n_1930),
		.B0(op_a[23]),
		.Y(n_1513));

	OAI21XL i_818557(
		.A0(n_1510),
		.A1(n_7350),
		.B0(n_6894),
		.Y(result[22]));

	AOI211X1 i_1315(
		.A0(n_1499),
		.A1(n_2293),
		.B0(n_6909),
		.C0(n_2311),
		.Y(n_1510));

	OAI21XL i_232(
		.A0(n_2303),
		.A1(n_1594),
		.B0(n_1496),
		.Y(n_1501));

	XNOR2X1 i_233(
		.A(op_a[22]),
		.B(n_2305),
		.Y(n_1500));

	OAI2BB1X1 i_234(
		.A0N(n_1587),
		.A1N(n_7326),
		.B0(n_7344),
		.Y(n_1499));

	NOR2X1 i_221376(
		.A(op_b[22]),
		.B(op_a[22]),
		.Y(n_1497));

	NAND2X1 i_1273(
		.A(n_1594),
		.B(n_2303),
		.Y(n_1496));

	AOI211X1 i_352(
		.A0(n_2198),
		.A1(n_2234),
		.B0(n_2233),
		.C0(n_1493),
		.Y(n_1494));

	NOR4BX1 i_1267(
		.AN(n_2234),
		.B(n_1339),
		.C(n_1297),
		.D(n_1392),
		.Y(n_1493));

	NOR2X1 i_211375(
		.A(op_b[21]),
		.B(op_a[21]),
		.Y(n_1492));

	OAI211X1 i_435(
		.A0(n_2229),
		.A1(n_2193),
		.B0(n_2228),
		.C0(n_1486),
		.Y(n_1487));

	NAND4BXL i_1257(
		.AN(n_2194),
		.B(n_1383),
		.C(n_929),
		.D(n_1385),
		.Y(n_1486));

	NAND2BX1 i_537100(
		.AN(op_a[21]),
		.B(op_b[21]),
		.Y(n_1485));

	OAI21XL i_828558(
		.A0(n_1482),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[21]));

	AOI211X1 i_1306(
		.A0(n_1471),
		.A1(n_2276),
		.B0(n_7335),
		.C0(n_2291),
		.Y(n_1482));

	OAI21XL i_225(
		.A0(n_2282),
		.A1(n_1567),
		.B0(n_1469),
		.Y(n_1473));

	AOI21X1 i_226(
		.A0(op_a[21]),
		.A1(n_2285),
		.B0(n_1464),
		.Y(n_1472));

	OAI2BB1X1 i_228(
		.A0N(n_1561),
		.A1N(n_7326),
		.B0(n_1716),
		.Y(n_1471));

	NAND2X1 i_1233(
		.A(n_1567),
		.B(n_2282),
		.Y(n_1469));

	AOI211X1 i_351(
		.A0(n_1843),
		.A1(n_1877),
		.B0(n_1838),
		.C0(n_1466),
		.Y(n_1467));

	NOR4BX1 i_1228(
		.AN(n_1877),
		.B(n_1297),
		.C(n_1293),
		.D(n_1365),
		.Y(n_1466));

	NOR2X1 i_1226(
		.A(n_2285),
		.B(op_a[21]),
		.Y(n_1464));

	OAI211X1 i_434(
		.A0(n_1804),
		.A1(n_1770),
		.B0(n_1765),
		.C0(n_1461),
		.Y(n_1462));

	NAND4BXL i_1218(
		.AN(n_1804),
		.B(n_1360),
		.C(n_931),
		.D(n_1286),
		.Y(n_1461));

	OAI21XL i_838559(
		.A0(n_1459),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[20]));

	AOI211X1 i_1297(
		.A0(n_1448),
		.A1(n_2258),
		.B0(n_7335),
		.C0(n_2274),
		.Y(n_1459));

	OAI21XL i_217(
		.A0(n_2268),
		.A1(n_1541),
		.B0(n_1445),
		.Y(n_1450));

	XNOR2X1 i_218(
		.A(op_a[20]),
		.B(n_1903),
		.Y(n_1449));

	OAI2BB1X1 i_219(
		.A0N(n_1534),
		.A1N(n_3062),
		.B0(n_1716),
		.Y(n_1448));

	NOR2X1 i_201374(
		.A(op_b[20]),
		.B(op_a[20]),
		.Y(n_1446));

	NAND2X1 i_1195(
		.A(n_1541),
		.B(n_2268),
		.Y(n_1445));

	AOI211X1 i_350(
		.A0(n_2167),
		.A1(n_2199),
		.B0(n_2198),
		.C0(n_1442),
		.Y(n_1443));

	NOR4BX1 i_1190(
		.AN(n_2168),
		.B(n_1339),
		.C(n_1297),
		.D(n_1340),
		.Y(n_1442));

	NOR2X1 i_191373(
		.A(op_b[19]),
		.B(op_a[19]),
		.Y(n_1441));

	OAI211X1 i_433(
		.A0(n_2162),
		.A1(n_2194),
		.B0(n_2193),
		.C0(n_1435),
		.Y(n_1436));

	NAND4BXL i_1181(
		.AN(n_2194),
		.B(n_1286),
		.C(n_1334),
		.D(n_933),
		.Y(n_1435));

	NAND2BX1 i_517098(
		.AN(op_a[19]),
		.B(op_b[19]),
		.Y(n_1434));

	OAI21XL i_848560(
		.A0(n_1431),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[19]));

	AOI211X1 i_1288(
		.A0(n_1420),
		.A1(n_2248),
		.B0(n_7335),
		.C0(n_2256),
		.Y(n_1431));

	OAI21XL i_167(
		.A0(n_2250),
		.A1(n_906),
		.B0(n_1418),
		.Y(n_1422));

	AOI21X1 i_186(
		.A0(op_a[19]),
		.A1(n_1930),
		.B0(n_1413),
		.Y(n_1421));

	OAI2BB1X1 i_188(
		.A0N(n_946),
		.A1N(n_3062),
		.B0(n_1716),
		.Y(n_1420));

	NAND2X1 i_1157(
		.A(n_906),
		.B(n_2250),
		.Y(n_1418));

	AOI211X1 i_348(
		.A0(n_1846),
		.A1(n_1847),
		.B0(n_1843),
		.C0(n_1415),
		.Y(n_1416));

	NOR4BX1 i_1151(
		.AN(n_1875),
		.B(n_1297),
		.C(n_1293),
		.D(n_903),
		.Y(n_1415));

	NOR2X1 i_1149(
		.A(n_1930),
		.B(op_a[19]),
		.Y(n_1413));

	OAI211X1 i_432(
		.A0(n_1773),
		.A1(n_1774),
		.B0(n_1770),
		.C0(n_1410),
		.Y(n_1411));

	NAND4BXL i_1143(
		.AN(n_1802),
		.B(n_931),
		.C(n_1286),
		.D(n_943),
		.Y(n_1410));

	OAI21XL i_858561(
		.A0(n_1408),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[18]));

	AOI211X1 i_1279(
		.A0(n_1397),
		.A1(n_2227),
		.B0(n_7335),
		.C0(n_2246),
		.Y(n_1408));

	OAI21XL i_130(
		.A0(n_2237),
		.A1(n_1494),
		.B0(n_1394),
		.Y(n_1399));

	AOI31X1 i_131(
		.A0(n_2174),
		.A1(op_a[18]),
		.A2(n_2239),
		.B0(n_1387),
		.Y(n_1398));

	OAI2BB1X1 i_132(
		.A0N(n_1487),
		.A1N(n_3062),
		.B0(n_1716),
		.Y(n_1397));

	NOR2X1 i_181372(
		.A(op_b[18]),
		.B(op_a[18]),
		.Y(n_1395));

	NAND2X1 i_1121(
		.A(n_1494),
		.B(n_2237),
		.Y(n_1394));

	AOI211X1 i_347(
		.A0(n_2132),
		.A1(n_2168),
		.B0(n_2167),
		.C0(n_1391),
		.Y(n_1392));

	NOR4BX1 i_1115(
		.AN(n_2168),
		.B(n_1244),
		.C(n_1198),
		.D(n_1294),
		.Y(n_1391));

	NOR2X1 i_171371(
		.A(op_b[17]),
		.B(op_a[17]),
		.Y(n_1390));

	AOI21X1 i_1112(
		.A0(n_2239),
		.A1(n_2174),
		.B0(op_a[18]),
		.Y(n_1387));

	OAI211X1 i_431(
		.A0(n_2163),
		.A1(n_2127),
		.B0(n_2162),
		.C0(n_1384),
		.Y(n_1385));

	NAND4BXL i_1105(
		.AN(n_2128),
		.B(n_1286),
		.C(n_933),
		.D(n_1287),
		.Y(n_1384));

	NAND2BX1 i_497096(
		.AN(op_a[17]),
		.B(op_b[17]),
		.Y(n_1383));

	OAI21XL i_868562(
		.A0(n_1380),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[17]));

	AOI211X1 i_1270(
		.A0(n_1369),
		.A1(n_2210),
		.B0(n_7335),
		.C0(n_2225),
		.Y(n_1380));

	OAI21XL i_125(
		.A0(n_2216),
		.A1(n_1467),
		.B0(n_1367),
		.Y(n_1371));

	AOI31X1 i_126(
		.A0(n_2153),
		.A1(op_a[17]),
		.A2(n_2218),
		.B0(n_1362),
		.Y(n_1370));

	OAI2BB1X1 i_127(
		.A0N(n_1462),
		.A1N(n_3062),
		.B0(n_1716),
		.Y(n_1369));

	NAND2X1 i_1075(
		.A(n_1467),
		.B(n_2216),
		.Y(n_1367));

	AOI211X1 i_346(
		.A0(n_1851),
		.A1(n_1875),
		.B0(n_1846),
		.C0(n_1364),
		.Y(n_1365));

	NOR4BX1 i_1070(
		.AN(n_1875),
		.B(n_1198),
		.C(n_1193),
		.D(n_1268),
		.Y(n_1364));

	AOI21X1 i_1068(
		.A0(n_2218),
		.A1(n_2153),
		.B0(op_a[17]),
		.Y(n_1362));

	OAI211X1 i_430(
		.A0(n_1802),
		.A1(n_1778),
		.B0(n_1773),
		.C0(n_1359),
		.Y(n_1360));

	NAND4BXL i_1061(
		.AN(n_1802),
		.B(n_1264),
		.C(n_935),
		.D(n_1186),
		.Y(n_1359));

	OAI21XL i_878563(
		.A0(n_1357),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[16]));

	AOI211X1 i_1261(
		.A0(n_1346),
		.A1(n_2192),
		.B0(n_7335),
		.C0(n_2208),
		.Y(n_1357));

	OAI21XL i_120(
		.A0(n_2202),
		.A1(n_1443),
		.B0(n_1343),
		.Y(n_1348));

	AOI21X1 i_121(
		.A0(op_a[16]),
		.A1(n_1899),
		.B0(n_1337),
		.Y(n_1347));

	OAI2BB1X1 i_122(
		.A0N(n_1436),
		.A1N(n_3062),
		.B0(n_1716),
		.Y(n_1346));

	NOR2X1 i_161370(
		.A(op_b[16]),
		.B(op_a[16]),
		.Y(n_1344));

	NAND2X1 i_1041(
		.A(n_1443),
		.B(n_2202),
		.Y(n_1343));

	NOR4BX1 i_345(
		.AN(n_2103),
		.B(n_1244),
		.C(n_1198),
		.D(n_1245),
		.Y(n_1341));

	AOI211X1 i_1038(
		.A0(n_2102),
		.A1(n_2133),
		.B0(n_2132),
		.C0(n_1341),
		.Y(n_1340));

	NOR2X1 i_151369(
		.A(op_b[15]),
		.B(op_a[15]),
		.Y(n_1339));

	NOR2X1 i_1035(
		.A(n_1899),
		.B(op_a[16]),
		.Y(n_1337));

	OAI211X1 i_429(
		.A0(n_2097),
		.A1(n_2128),
		.B0(n_2127),
		.C0(n_1333),
		.Y(n_1334));

	NAND4BXL i_1029(
		.AN(n_2128),
		.B(n_1186),
		.C(n_1238),
		.D(n_937),
		.Y(n_1333));

	NAND2BX1 i_477094(
		.AN(op_a[15]),
		.B(op_b[15]),
		.Y(n_1332));

	OAI21XL i_888564(
		.A0(n_1329),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[15]));

	AOI211X1 i_1252(
		.A0(n_1318),
		.A1(n_2182),
		.B0(n_6909),
		.C0(n_2190),
		.Y(n_1329));

	OAI21XL i_115(
		.A0(n_2184),
		.A1(n_1416),
		.B0(n_1316),
		.Y(n_1320));

	AOI31X1 i_116(
		.A0(n_1924),
		.A1(op_a[15]),
		.A2(n_1926),
		.B0(n_1314),
		.Y(n_1319));

	OAI2BB1X1 i_117(
		.A0N(n_1411),
		.A1N(n_7326),
		.B0(n_1716),
		.Y(n_1318));

	NAND2X1 i_1008(
		.A(n_1416),
		.B(n_2184),
		.Y(n_1316));

	AOI21X1 i_1006(
		.A0(n_1926),
		.A1(n_1924),
		.B0(op_a[15]),
		.Y(n_1314));

	OAI21XL i_898565(
		.A0(n_1310),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[14]));

	AOI211X1 i_1243(
		.A0(n_1299),
		.A1(n_2161),
		.B0(n_6909),
		.C0(n_2180),
		.Y(n_1310));

	OAI21XL i_110(
		.A0(n_2171),
		.A1(n_1392),
		.B0(n_1296),
		.Y(n_1301));

	AOI21X1 i_111(
		.A0(n_7270),
		.A1(n_2174),
		.B0(n_1291),
		.Y(n_1300));

	OAI2BB1X1 i_112(
		.A0N(n_1385),
		.A1N(n_7326),
		.B0(n_1716),
		.Y(n_1299));

	NOR2X1 i_141368(
		.A(op_b[14]),
		.B(op_a[14]),
		.Y(n_1297));

	NAND2X1 i_984(
		.A(n_1392),
		.B(n_2171),
		.Y(n_1296));

	AOI211X1 i_981(
		.A0(n_2066),
		.A1(n_2103),
		.B0(n_2102),
		.C0(n_855),
		.Y(n_1294));

	NOR2X1 i_131367(
		.A(op_b[13]),
		.B(op_a[13]),
		.Y(n_1293));

	NOR2X1 i_978(
		.A(n_2174),
		.B(n_7270),
		.Y(n_1291));

	NAND4X1 i_426(
		.A(n_1186),
		.B(n_937),
		.C(n_1187),
		.D(n_2062),
		.Y(n_1288));

	OAI211X1 i_972(
		.A0(n_2098),
		.A1(n_2061),
		.B0(n_2097),
		.C0(n_1288),
		.Y(n_1287));

	NAND2BX1 i_457092(
		.AN(op_a[13]),
		.B(op_b[13]),
		.Y(n_1286));

	OAI21XL i_908566(
		.A0(n_1283),
		.A1(n_7347),
		.B0(n_6894),
		.Y(result[13]));

	AOI211X1 i_1234(
		.A0(n_1272),
		.A1(n_2144),
		.B0(n_6909),
		.C0(n_2159),
		.Y(n_1283));

	OAI21XL i_105(
		.A0(n_2150),
		.A1(n_1365),
		.B0(n_1270),
		.Y(n_1274));

	AOI21X1 i_106(
		.A0(op_a[13]),
		.A1(n_2153),
		.B0(n_1267),
		.Y(n_1273));

	OAI2BB1X1 i_107(
		.A0N(n_1360),
		.A1N(n_7326),
		.B0(n_1716),
		.Y(n_1272));

	NAND2X1 i_950(
		.A(n_1365),
		.B(n_2150),
		.Y(n_1270));

	AOI31X1 i_947(
		.A0(n_1873),
		.A1(n_1863),
		.A2(n_1167),
		.B0(n_3092),
		.Y(n_1268));

	NOR2X1 i_945(
		.A(n_2153),
		.B(op_a[13]),
		.Y(n_1267));

	OAI31X1 i_939(
		.A0(n_1800),
		.A1(n_1790),
		.A2(n_1162),
		.B0(n_2080),
		.Y(n_1264));

	OAI21XL i_918567(
		.A0(n_1262),
		.A1(n_7347),
		.B0(n_6893),
		.Y(result[12]));

	AOI211X1 i_1225(
		.A0(n_1251),
		.A1(n_2126),
		.B0(n_6909),
		.C0(n_2142),
		.Y(n_1262));

	OAI21XL i_99(
		.A0(n_2136),
		.A1(n_1340),
		.B0(n_1248),
		.Y(n_1253));

	XNOR2X1 i_100(
		.A(n_1895),
		.B(op_a[12]),
		.Y(n_1252));

	OAI2BB1X1 i_101(
		.A0N(n_1334),
		.A1N(n_7326),
		.B0(n_7344),
		.Y(n_1251));

	NOR2X1 i_121366(
		.A(op_b[12]),
		.B(op_a[12]),
		.Y(n_1249));

	NAND2X1 i_918(
		.A(n_1340),
		.B(n_2136),
		.Y(n_1248));

	NOR4BX1 i_336(
		.AN(n_2039),
		.B(n_1144),
		.C(n_1100),
		.D(n_2004),
		.Y(n_1246));

	AOI211X1 i_915(
		.A0(n_2038),
		.A1(n_2067),
		.B0(n_2066),
		.C0(n_1246),
		.Y(n_1245));

	NOR2X1 i_111365(
		.A(op_b[11]),
		.B(op_a[11]),
		.Y(n_1244));

	NAND4X1 i_422(
		.A(n_1090),
		.B(n_2062),
		.C(n_1137),
		.D(n_942),
		.Y(n_1239));

	NAND3X1 i_908(
		.A(n_2061),
		.B(n_1239),
		.C(n_862),
		.Y(n_1238));

	NAND2BX1 i_437090(
		.AN(op_a[11]),
		.B(op_b[11]),
		.Y(n_1237));

	OAI21XL i_928568(
		.A0(n_1234),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[11]));

	AOI211X1 i_1216(
		.A0(n_1223),
		.A1(n_2116),
		.B0(n_6909),
		.C0(n_2124),
		.Y(n_1234));

	OAI21XL i_94(
		.A0(n_2118),
		.A1(n_903),
		.B0(n_1221),
		.Y(n_1225));

	AOI21X1 i_95(
		.A0(op_a[11]),
		.A1(n_1924),
		.B0(n_1217),
		.Y(n_1224));

	OAI2BB1X1 i_96(
		.A0N(n_943),
		.A1N(n_7326),
		.B0(n_7344),
		.Y(n_1223));

	NAND2X1 i_886(
		.A(n_903),
		.B(n_2118),
		.Y(n_1221));

	NOR4BX1 i_334(
		.AN(n_1863),
		.B(n_1053),
		.C(n_1097),
		.D(n_1870),
		.Y(n_1219));

	AOI211X1 i_883(
		.A0(n_1862),
		.A1(n_1863),
		.B0(n_1859),
		.C0(n_1219),
		.Y(n_1218));

	NOR2X1 i_881(
		.A(n_1924),
		.B(op_a[11]),
		.Y(n_1217));

	AOI211X1 i_877(
		.A0(n_1797),
		.A1(n_1799),
		.B0(n_861),
		.C0(n_1786),
		.Y(n_1213));

	OAI21XL i_938569(
		.A0(n_1211),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[10]));

	AOI211X1 i_1207(
		.A0(n_1200),
		.A1(n_2096),
		.B0(n_6909),
		.C0(n_2114),
		.Y(n_1211));

	OAI21XL i_89(
		.A0(n_2106),
		.A1(n_1294),
		.B0(n_1197),
		.Y(n_1202));

	AOI21X1 i_90(
		.A0(n_7290),
		.A1(n_2108),
		.B0(n_1191),
		.Y(n_1201));

	OAI2BB1X1 i_91(
		.A0N(n_1287),
		.A1N(n_7326),
		.B0(n_7344),
		.Y(n_1200));

	NOR2X1 i_101364(
		.A(op_b[10]),
		.B(op_a[10]),
		.Y(n_1198));

	NAND2X1 i_856(
		.A(n_1294),
		.B(n_2106),
		.Y(n_1197));

	AOI31X1 i_853(
		.A0(n_2039),
		.A1(n_2003),
		.A2(n_1976),
		.B0(n_3089),
		.Y(n_1194));

	NOR2X1 i_91363(
		.A(op_b[9]),
		.B(op_a[9]),
		.Y(n_1193));

	NOR2X1 i_851(
		.A(n_2108),
		.B(n_7290),
		.Y(n_1191));

	NAND4BXL i_418(
		.AN(n_1997),
		.B(n_1090),
		.C(n_942),
		.D(n_1972),
		.Y(n_1188));

	NAND4X1 i_846(
		.A(n_1089),
		.B(n_1785),
		.C(n_1188),
		.D(n_860),
		.Y(n_1187));

	NAND2BX1 i_417088(
		.AN(op_a[9]),
		.B(op_b[9]),
		.Y(n_1186));

	OAI21XL i_948570(
		.A0(n_1183),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[9]));

	AOI211X1 i_1198(
		.A0(n_1172),
		.A1(n_2079),
		.B0(n_6909),
		.C0(n_2094),
		.Y(n_1183));

	OAI21XL i_84(
		.A0(n_2085),
		.A1(n_1268),
		.B0(n_1170),
		.Y(n_1174));

	AOI31X1 i_85(
		.A0(n_2017),
		.A1(op_a[9]),
		.A2(n_2087),
		.B0(n_1166),
		.Y(n_1173));

	OAI2BB1X1 i_86(
		.A0N(n_1264),
		.A1N(n_7326),
		.B0(n_7344),
		.Y(n_1172));

	NAND2X1 i_824(
		.A(n_1268),
		.B(n_2085),
		.Y(n_1170));

	NAND3X1 i_18(
		.A(n_1869),
		.B(n_3085),
		.C(n_1871),
		.Y(n_1168));

	NAND2X1 i_821(
		.A(n_1168),
		.B(n_2020),
		.Y(n_1167));

	AOI21X1 i_820(
		.A0(n_2087),
		.A1(n_2017),
		.B0(op_a[9]),
		.Y(n_1166));

	AOI2BB1X1 i_814(
		.A0N(n_1798),
		.A1N(n_857),
		.B0(n_2013),
		.Y(n_1162));

	OAI21XL i_958571(
		.A0(n_1160),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[8]));

	AOI211X1 i_1189(
		.A0(n_1149),
		.A1(n_2060),
		.B0(n_6909),
		.C0(n_2077),
		.Y(n_1160));

	OAI21XL i_79(
		.A0(n_2070),
		.A1(n_1245),
		.B0(n_1146),
		.Y(n_1151));

	XNOR2X1 i_80(
		.A(op_a[8]),
		.B(n_1891),
		.Y(n_1150));

	OAI2BB1X1 i_81(
		.A0N(n_1238),
		.A1N(n_7326),
		.B0(n_7344),
		.Y(n_1149));

	NOR2X1 i_81362(
		.A(op_b[8]),
		.B(op_a[8]),
		.Y(n_1147));

	NAND2X1 i_794(
		.A(n_1245),
		.B(n_2070),
		.Y(n_1146));

	NOR2X1 i_7(
		.A(op_b[7]),
		.B(op_a[7]),
		.Y(n_1144));

	OAI21XL i_784(
		.A0(n_856),
		.A1(n_1997),
		.B0(n_1998),
		.Y(n_1137));

	NOR2BX1 i_337080(
		.AN(op_b[1]),
		.B(op_a[1]),
		.Y(n_1136));

	NAND2BX1 i_397086(
		.AN(op_a[7]),
		.B(op_b[7]),
		.Y(n_1135));

	OAI21XL i_968572(
		.A0(n_1132),
		.A1(n_7347),
		.B0(n_6893),
		.Y(result[7]));

	AOI21X1 i_1180(
		.A0(n_1122),
		.A1(n_2049),
		.B0(n_2059),
		.Y(n_1132));

	AOI21X1 i_768(
		.A0(n_1915),
		.A1(n_2052),
		.B0(n_1917),
		.Y(n_1129));

	OAI21XL i_73(
		.A0(n_2053),
		.A1(n_1218),
		.B0(n_1119),
		.Y(n_1123));

	OAI2BB1X1 i_74(
		.A0N(n_3076),
		.A1N(n_7369),
		.B0(n_7329),
		.Y(n_1122));

	NAND2X1 i_763(
		.A(n_1218),
		.B(n_2053),
		.Y(n_1119));

	NOR2X1 i_759(
		.A(op_a[7]),
		.B(n_2051),
		.Y(n_1116));

	OAI21XL i_978573(
		.A0(n_1113),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[6]));

	AOI21X1 i_1171(
		.A0(n_1103),
		.A1(n_2028),
		.B0(n_2048),
		.Y(n_1113));

	AOI21X1 i_744(
		.A0(n_1915),
		.A1(n_2037),
		.B0(n_1917),
		.Y(n_1110));

	OAI21XL i_66(
		.A0(n_2042),
		.A1(n_1194),
		.B0(n_1099),
		.Y(n_1104));

	OAI2BB1X1 i_67(
		.A0N(n_1187),
		.A1N(n_3062),
		.B0(n_7329),
		.Y(n_1103));

	NOR2X1 i_61361(
		.A(op_b[6]),
		.B(op_a[6]),
		.Y(n_1100));

	NAND2X1 i_739(
		.A(n_1194),
		.B(n_2042),
		.Y(n_1099));

	NOR2X1 i_31360(
		.A(op_b[3]),
		.B(op_a[3]),
		.Y(n_1097));

	NOR2X1 i_21359(
		.A(op_b[2]),
		.B(op_a[2]),
		.Y(n_1096));

	NOR2X1 i_5(
		.A(op_b[5]),
		.B(op_a[5]),
		.Y(n_1095));

	NOR2X1 i_732(
		.A(op_a[6]),
		.B(n_2036),
		.Y(n_1092));

	NAND2BX1 i_377084(
		.AN(op_a[5]),
		.B(op_b[5]),
		.Y(n_1090));

	NAND2X1 i_726(
		.A(n_1090),
		.B(n_1787),
		.Y(n_1089));

	OAI21XL i_988574(
		.A0(n_1087),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[5]));

	NOR4BX1 i_1162(
		.AN(n_1085),
		.B(n_1084),
		.C(n_2025),
		.D(n_1076),
		.Y(n_1087));

	NAND4X1 i_715(
		.A(n_1785),
		.B(n_1090),
		.C(n_1162),
		.D(n_3062),
		.Y(n_1085));

	AOI21X1 i_712(
		.A0(n_1915),
		.A1(n_2019),
		.B0(n_1917),
		.Y(n_1084));

	AOI31X1 i_60(
		.A0(n_1168),
		.A1(n_2020),
		.A2(n_2021),
		.B0(n_1073),
		.Y(n_1078));

	AOI22X1 i_713(
		.A0(n_7344),
		.A1(n_1071),
		.B0(n_1785),
		.B1(n_1090),
		.Y(n_1076));

	AOI21X1 i_706(
		.A0(n_1168),
		.A1(n_2020),
		.B0(n_2021),
		.Y(n_1073));

	NOR2X1 i_1(
		.A(op_b[1]),
		.B(op_a[1]),
		.Y(n_1072));

	NAND2BX1 i_703(
		.AN(n_1162),
		.B(n_3062),
		.Y(n_1071));

	NOR2X1 i_701(
		.A(op_a[5]),
		.B(n_2018),
		.Y(n_1070));

	NAND2BX1 i_347081(
		.AN(op_a[2]),
		.B(op_b[2]),
		.Y(n_1068));

	OAI21XL i_998575(
		.A0(n_1066),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[4]));

	AOI21X1 i_1153(
		.A0(n_1056),
		.A1(n_1995),
		.B0(n_2011),
		.Y(n_1066));

	AOI21X1 i_681(
		.A0(n_1915),
		.A1(n_2001),
		.B0(n_1917),
		.Y(n_1063));

	OAI21XL i_55(
		.A0(n_2005),
		.A1(n_2004),
		.B0(n_1052),
		.Y(n_1057));

	OAI2BB1X1 i_56(
		.A0N(n_1137),
		.A1N(n_3062),
		.B0(n_7329),
		.Y(n_1056));

	NOR2X1 i_4(
		.A(op_b[4]),
		.B(op_a[4]),
		.Y(n_1053));

	NAND2X1 i_676(
		.A(n_2004),
		.B(n_2005),
		.Y(n_1052));

	NOR2X1 i_670(
		.A(op_a[4]),
		.B(n_2000),
		.Y(n_1048));

	NAND2BX1 i_357082(
		.AN(n_7302),
		.B(op_b[3]),
		.Y(n_1045));

	OAI21XL i_1008576(
		.A0(n_1042),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[3]));

	AOI21X1 i_1144(
		.A0(n_1032),
		.A1(n_1984),
		.B0(n_1994),
		.Y(n_1042));

	AOI21X1 i_651(
		.A0(n_1915),
		.A1(n_1987),
		.B0(n_1917),
		.Y(n_1039));

	OAI21XL i_49(
		.A0(n_1988),
		.A1(n_1870),
		.B0(n_1029),
		.Y(n_1033));

	OAI2BB1X1 i_50(
		.A0N(n_1797),
		.A1N(n_7369),
		.B0(n_7329),
		.Y(n_1032));

	NAND2X1 i_646(
		.A(n_1870),
		.B(n_1988),
		.Y(n_1029));

	NOR2X1 i_642(
		.A(n_7302),
		.B(n_1986),
		.Y(n_1026));

	OAI21XL i_1018577(
		.A0(n_1023),
		.A1(n_7350),
		.B0(n_6893),
		.Y(result[2]));

	AOI21X1 i_1135(
		.A0(n_1013),
		.A1(n_1970),
		.B0(n_1983),
		.Y(n_1023));

	AOI21X1 i_627(
		.A0(n_1915),
		.A1(n_1975),
		.B0(n_1917),
		.Y(n_1020));

	XOR2X1 i_43(
		.A(n_1976),
		.B(n_1977),
		.Y(n_1014));

	OAI2BB1X1 i_44(
		.A0N(n_1972),
		.A1N(n_7369),
		.B0(n_7329),
		.Y(n_1013));

	NOR2X1 i_617(
		.A(op_a[2]),
		.B(n_1974),
		.Y(n_1006));

	OAI21XL i_1028578(
		.A0(n_1002),
		.A1(n_7350),
		.B0(n_6893),
		.Y(result[1]));

	AOI21X1 i_1126(
		.A0(n_992),
		.A1(n_1959),
		.B0(n_1969),
		.Y(n_1002));

	AOI21X1 i_601(
		.A0(n_1915),
		.A1(n_1962),
		.B0(n_1917),
		.Y(n_999));

	OAI31X1 i_37(
		.A0(n_3083),
		.A1(n_1072),
		.A2(n_3085),
		.B0(n_988),
		.Y(n_993));

	OAI2BB1X1 i_38(
		.A0N(n_1795),
		.A1N(n_7369),
		.B0(n_7329),
		.Y(n_992));

	OAI21XL i_595(
		.A0(n_1072),
		.A1(n_3083),
		.B0(n_3085),
		.Y(n_988));

	NOR2X1 i_592(
		.A(op_a[1]),
		.B(n_1961),
		.Y(n_986));

	AOI21X1 i_1038579(
		.A0(n_983),
		.A1(n_9076575),
		.B0(n_827),
		.Y(n_984));

	NAND3BX1 i_1117(
		.AN(n_981),
		.B(n_1957),
		.C(n_976),
		.Y(n_983));

	AOI21X1 i_582(
		.A0(n_7344),
		.A1(n_6939),
		.B0(n_1795),
		.Y(n_981));

	OR2X1 i_34(
		.A(n_1946),
		.B(n_974),
		.Y(n_978));

	OAI21XL i_583(
		.A0(n_973),
		.A1(n_1955),
		.B0(op_a[0]),
		.Y(n_976));

	NOR2X1 i_574(
		.A(n_3085),
		.B(n_3095),
		.Y(n_974));

	AOI21X1 i_575(
		.A0(n_7344),
		.A1(n_7323),
		.B0(op_b[0]),
		.Y(n_973));

	NOR3X1 i_570(
		.A(n_1950),
		.B(op_a[31]),
		.C(n_1733),
		.Y(n_971));

	NOR2X1 i_569(
		.A(op_b[31]),
		.B(n_3095),
		.Y(n_970));

	NAND4X1 i_559(
		.A(n_1936),
		.B(n_1915),
		.C(n_1938),
		.D(n_1918),
		.Y(n_967));

	AOI22X1 i_291(
		.A0(n_1810),
		.A1(n_3062),
		.B0(n_1883),
		.B1(n_6904),
		.Y(n_964));

	NAND3X1 i_292(
		.A(n_958),
		.B(n_1944),
		.C(n_6901),
		.Y(n_963));

	OAI221XL i_293(
		.A0(n_3095),
		.A1(n_1883),
		.B0(n_1810),
		.B1(n_1738),
		.C0(n_1716),
		.Y(n_962));

	NAND2X1 i_550(
		.A(cmd[1]),
		.B(op_b[31]),
		.Y(n_958));

	OAI21XL i_452(
		.A0(n_951),
		.A1(n_1713),
		.B0(n_885),
		.Y(n_955));

	NAND2BX1 i_455(
		.AN(op_a[30]),
		.B(op_b[30]),
		.Y(n_954));

	NOR2BX1 i_542(
		.AN(op_a[30]),
		.B(op_b[30]),
		.Y(n_952));

	AOI2BB1X1 i_453(
		.A0N(n_949),
		.A1N(n_1743),
		.B0(n_3070),
		.Y(n_951));

	AOI21X1 i_454(
		.A0(n_1612),
		.A1(n_1809),
		.B0(n_1751),
		.Y(n_949));

	OAI211X1 i_436(
		.A0(n_1765),
		.A1(n_1766),
		.B0(n_1762),
		.C0(n_945),
		.Y(n_946));

	NAND4BXL i_535(
		.AN(n_1804),
		.B(n_927),
		.C(n_1383),
		.D(n_1411),
		.Y(n_945));

	OR3XL i_428(
		.A(n_1782),
		.B(n_1800),
		.C(n_1213),
		.Y(n_944));

	OAI211X1 i_533(
		.A0(n_1781),
		.A1(n_1782),
		.B0(n_1778),
		.C0(n_944),
		.Y(n_943));

	NAND2BX1 i_367083(
		.AN(op_a[4]),
		.B(op_b[4]),
		.Y(n_942));

	NOR2BX1 i_387085(
		.AN(op_b[6]),
		.B(op_a[6]),
		.Y(n_940));

	NAND2BX1 i_407087(
		.AN(op_a[8]),
		.B(op_b[8]),
		.Y(n_937));

	NAND2BX1 i_427089(
		.AN(n_7290),
		.B(op_b[10]),
		.Y(n_935));

	NAND2BX1 i_447091(
		.AN(op_a[12]),
		.B(op_b[12]),
		.Y(n_933));

	NAND2BX1 i_467093(
		.AN(n_7270),
		.B(op_b[14]),
		.Y(n_931));

	NAND2BX1 i_487095(
		.AN(op_a[16]),
		.B(op_b[16]),
		.Y(n_929));

	NAND2BX1 i_507097(
		.AN(op_a[18]),
		.B(op_b[18]),
		.Y(n_927));

	NAND2BX1 i_527099(
		.AN(op_a[20]),
		.B(op_b[20]),
		.Y(n_925));

	NAND2BX1 i_547101(
		.AN(op_a[22]),
		.B(op_b[22]),
		.Y(n_923));

	NAND2BX1 i_567103(
		.AN(op_a[24]),
		.B(op_b[24]),
		.Y(n_921));

	OAI21XL i_367(
		.A0(n_913),
		.A1(n_1703),
		.B0(n_1812),
		.Y(n_917));

	OAI21XL i_514(
		.A0(op_a[30]),
		.A1(op_b[30]),
		.B0(n_917),
		.Y(n_915));

	AOI21X1 i_368(
		.A0(n_1816),
		.A1(n_3086),
		.B0(n_1815),
		.Y(n_913));

	AOI211X1 i_369(
		.A0(n_1822),
		.A1(n_1823),
		.B0(n_1819),
		.C0(n_909),
		.Y(n_911));

	NOR2X1 i_510(
		.A(n_1617),
		.B(n_1882),
		.Y(n_909));

	AOI211X1 i_353(
		.A0(n_1838),
		.A1(n_1839),
		.B0(n_1835),
		.C0(n_905),
		.Y(n_906));

	NOR4BX1 i_506(
		.AN(n_1877),
		.B(n_1395),
		.C(n_1390),
		.D(n_1416),
		.Y(n_905));

	NOR4BX1 i_342(
		.AN(n_1873),
		.B(n_1198),
		.C(n_1193),
		.D(n_1218),
		.Y(n_904));

	AOI211X1 i_504(
		.A0(n_1854),
		.A1(n_1855),
		.B0(n_1851),
		.C0(n_904),
		.Y(n_903));

	NAND2BX1 i_937140(
		.AN(op_b[29]),
		.B(op_a[29]),
		.Y(n_885));

	NAND2BX1 i_412(
		.AN(n_2324),
		.B(n_2362),
		.Y(n_882));

	NAND2BX1 i_409(
		.AN(n_1757),
		.B(n_1758),
		.Y(n_879));

	NAND2X1 i_378(
		.A(n_2029),
		.B(n_2062),
		.Y(n_862));

	NOR2X1 i_377(
		.A(n_1789),
		.B(n_1790),
		.Y(n_861));

	NAND3X1 i_376(
		.A(n_1090),
		.B(n_942),
		.C(n_3087),
		.Y(n_860));

	NAND3X1 i_372(
		.A(n_1068),
		.B(n_1795),
		.C(n_3065),
		.Y(n_857));

	NAND2X1 i_371(
		.A(op_a[0]),
		.B(n_3065),
		.Y(n_856));

	NOR4BX1 i_332(
		.AN(n_2103),
		.B(n_1144),
		.C(n_1100),
		.D(n_1194),
		.Y(n_855));

	AOI31X1 i_33(
		.A0(op_a[31]),
		.A1(n_1733),
		.A2(n_1950),
		.B0(n_971),
		.Y(n_828));

	NOR2X1 i_9(
		.A(n_1733),
		.B(n_9076575),
		.Y(n_827));

	AOI22X1 i_1460(
		.A0(n_1613),
		.A1(n_7344),
		.B0(n_1640),
		.B1(n_3069),
		.Y(n_1620));

	AOI21X1 i_268(
		.A0(op_a[27]),
		.A1(n_1936),
		.B0(n_1614),
		.Y(n_1622));

	AOI21X1 i_267(
		.A0(n_2382),
		.A1(n_911),
		.B0(n_1618),
		.Y(n_1623));

	AND4X1 i_1463(
		.A(n_3069),
		.B(n_1640),
		.C(n_949),
		.D(n_3062),
		.Y(n_1630));

	NOR4X1 i_1360(
		.A(n_1630),
		.B(n_2387),
		.C(n_6909),
		.D(n_1620),
		.Y(n_1632));

	OAI21XL i_768552(
		.A0(n_1632),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[27]));

	NAND4BXL i_1476(
		.AN(n_2325),
		.B(n_1534),
		.C(n_1485),
		.D(n_925),
		.Y(n_1635));

	OAI211X1 i_448(
		.A0(n_2294),
		.A1(n_2325),
		.B0(n_2324),
		.C0(n_1635),
		.Y(n_1637));

	OAI2BB1X1 i_447(
		.A0N(n_1637),
		.A1N(n_2362),
		.B0(n_2361),
		.Y(n_1639));

	NAND2BX1 i_597106(
		.AN(op_a[27]),
		.B(op_b[27]),
		.Y(n_1640));

	NOR4BX1 i_1485(
		.AN(n_2300),
		.B(n_1539),
		.C(n_1497),
		.D(n_1541),
		.Y(n_1645));

	NOR2BX1 i_1487(
		.AN(n_2367),
		.B(n_1647),
		.Y(n_1646));

	AOI211X1 i_363(
		.A0(n_2299),
		.A1(n_2330),
		.B0(n_2329),
		.C0(n_1645),
		.Y(n_1647));

	OAI222XL i_1488(
		.A0(op_b[27]),
		.A1(op_a[27]),
		.B0(op_b[26]),
		.B1(op_a[26]),
		.C0(n_1646),
		.C1(n_2366),
		.Y(n_1648));

	NOR2X1 i_271381(
		.A(op_b[27]),
		.B(op_a[27]),
		.Y(n_1650));

	NAND2X1 i_1491(
		.A(n_2402),
		.B(n_2401),
		.Y(n_1652));

	NAND2BX1 i_1496(
		.AN(n_2390),
		.B(n_1654),
		.Y(n_1653));

	OAI21XL i_275(
		.A0(n_2393),
		.A1(n_7323),
		.B0(n_7344),
		.Y(n_1654));

	XNOR2X1 i_273(
		.A(op_a[28]),
		.B(n_1911),
		.Y(n_1655));

	OAI21XL i_272(
		.A0(n_2402),
		.A1(n_2401),
		.B0(n_1652),
		.Y(n_1656));

	NOR2X1 i_1497(
		.A(n_1655),
		.B(n_3068),
		.Y(n_1661));

	NAND4BXL i_1369(
		.AN(n_6909),
		.B(n_2397),
		.C(n_2404),
		.D(n_1653),
		.Y(n_1665));

	OAI2BB1X1 i_758551(
		.A0N(n_1665),
		.A1N(n_9076575),
		.B0(n_6894),
		.Y(result[28]));

	AOI31X1 i_449(
		.A0(n_1809),
		.A1(n_1758),
		.A2(n_1561),
		.B0(n_2408),
		.Y(n_1670));

	NOR2X1 i_1519(
		.A(n_2417),
		.B(op_a[29]),
		.Y(n_1672));

	NAND4BXL i_1522(
		.AN(n_1567),
		.B(n_1823),
		.C(n_1881),
		.D(n_1831),
		.Y(n_1674));

	AOI21X1 i_1525(
		.A0(n_1674),
		.A1(n_2411),
		.B0(n_3077),
		.Y(n_1676));

	OAI21XL i_1526(
		.A0(n_1676),
		.A1(n_1815),
		.B0(n_2413),
		.Y(n_1678));

	OAI2BB1X1 i_280(
		.A0N(n_2409),
		.A1N(n_7326),
		.B0(n_7344),
		.Y(n_1681));

	AOI21X1 i_279(
		.A0(op_a[29]),
		.A1(n_2417),
		.B0(n_1672),
		.Y(n_1682));

	OAI31X1 i_278(
		.A0(n_1676),
		.A1(n_1815),
		.A2(n_2413),
		.B0(n_1678),
		.Y(n_1683));

	NOR3X1 i_1535(
		.A(n_2409),
		.B(n_2406),
		.C(n_7323),
		.Y(n_1689));

	AOI211X1 i_1378(
		.A0(n_1681),
		.A1(n_2406),
		.B0(n_6909),
		.C0(n_2423),
		.Y(n_1692));

	OAI21XL i_748550(
		.A0(n_1692),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[29]));

	NOR4BX1 i_1554(
		.AN(n_2367),
		.B(n_1539),
		.C(n_1497),
		.D(n_1594),
		.Y(n_1696));

	NOR2X1 i_281382(
		.A(op_b[28]),
		.B(op_a[28]),
		.Y(n_1697));

	NOR3BX1 i_1557(
		.AN(n_1816),
		.B(n_1700),
		.C(n_1699),
		.Y(n_1698));

	AOI211X1 i_366(
		.A0(n_2329),
		.A1(n_2367),
		.B0(n_2366),
		.C0(n_1696),
		.Y(n_1699));

	NOR2X1 i_261380(
		.A(op_b[26]),
		.B(op_a[26]),
		.Y(n_1700));

	NOR2X1 i_291383(
		.A(op_b[29]),
		.B(op_a[29]),
		.Y(n_1703));

	AOI221X1 i_365(
		.A0(n_2399),
		.A1(n_3066),
		.B0(op_a[28]),
		.B1(op_b[28]),
		.C0(n_1698),
		.Y(n_1704));

	NAND3BX1 i_1561(
		.AN(n_2325),
		.B(n_2362),
		.C(n_1587),
		.Y(n_1705));

	NAND2BX1 i_607107(
		.AN(op_a[28]),
		.B(op_b[28]),
		.Y(n_1706));

	NAND3X1 i_451(
		.A(n_882),
		.B(n_2361),
		.C(n_1705),
		.Y(n_1708));

	NAND2BX1 i_587105(
		.AN(op_a[26]),
		.B(op_b[26]),
		.Y(n_1709));

	NOR2BX1 i_927139(
		.AN(op_a[28]),
		.B(op_b[28]),
		.Y(n_1710));

	NOR2BX1 i_617108(
		.AN(op_b[29]),
		.B(op_a[29]),
		.Y(n_1713));

	AOI221X1 i_450(
		.A0(n_2391),
		.A1(n_1706),
		.B0(n_1708),
		.B1(n_2426),
		.C0(n_1710),
		.Y(n_1714));

	NAND3BX1 i_1092(
		.AN(cmd[0]),
		.B(cmd[2]),
		.C(n_1736),
		.Y(n_1716));

	OAI21XL i_288(
		.A0(n_2434),
		.A1(n_6911),
		.B0(n_2436),
		.Y(n_1720));

	OAI221XL i_2879002(
		.A0(n_2431),
		.A1(n_3095),
		.B0(n_7323),
		.B1(n_3088),
		.C0(n_7344),
		.Y(n_1722));

	AOI22X1 i_285(
		.A0(n_3088),
		.A1(n_7326),
		.B0(n_2431),
		.B1(n_7341),
		.Y(n_1723));

	NOR2X1 i_10(
		.A(n_1915),
		.B(n_6911),
		.Y(n_1727));

	AOI21X1 i_1387(
		.A0(n_1722),
		.A1(n_2425),
		.B0(n_2441),
		.Y(n_1730));

	OAI21XL i_738549(
		.A0(n_1730),
		.A1(n_907),
		.B0(n_6893),
		.Y(result[30]));

	AOI21X1 i_1396(
		.A0(n_962),
		.A1(n_1740),
		.B0(n_1949),
		.Y(n_1733));

	NAND2X1 i_1587(
		.A(n_1733),
		.B(n_907),
		.Y(n_1734));

	OAI21XL i_728548(
		.A0(n_1733),
		.A1(n_907),
		.B0(n_1734),
		.Y(result[31]));

	NOR2X1 i_14(
		.A(cmd[3]),
		.B(cmd[1]),
		.Y(n_1736));

	NAND3BX1 i_1081(
		.AN(cmd[2]),
		.B(cmd[0]),
		.C(n_1736),
		.Y(n_1738));

	XOR2X1 i_1607206(
		.A(op_a[31]),
		.B(op_b[31]),
		.Y(n_1740));

	NOR2BX1 i_917138(
		.AN(op_a[27]),
		.B(op_b[27]),
		.Y(n_1741));

	AOI21X1 i_1897235(
		.A0(n_1706),
		.A1(n_1741),
		.B0(n_1710),
		.Y(n_1742));

	NAND2X1 i_13(
		.A(n_1706),
		.B(n_1640),
		.Y(n_1743));

	NOR2BX1 i_907137(
		.AN(op_a[26]),
		.B(op_b[26]),
		.Y(n_1744));

	NOR2BX1 i_897136(
		.AN(op_a[25]),
		.B(op_b[25]),
		.Y(n_1745));

	AOI21X1 i_1877233(
		.A0(n_1709),
		.A1(n_1745),
		.B0(n_1744),
		.Y(n_1746));

	NOR2BX1 i_887135(
		.AN(op_a[24]),
		.B(op_b[24]),
		.Y(n_1747));

	NOR2BX1 i_877134(
		.AN(op_a[23]),
		.B(op_b[23]),
		.Y(n_1748));

	AOI21X1 i_1857231(
		.A0(n_921),
		.A1(n_1748),
		.B0(n_1747),
		.Y(n_1749));

	NAND2X1 i_2197263(
		.A(n_1709),
		.B(n_1585),
		.Y(n_1750));

	OAI21XL i_2507290(
		.A0(n_1750),
		.A1(n_1749),
		.B0(n_1746),
		.Y(n_1751));

	NOR2BX1 i_867133(
		.AN(op_a[22]),
		.B(op_b[22]),
		.Y(n_1752));

	NOR2BX1 i_857132(
		.AN(op_a[21]),
		.B(op_b[21]),
		.Y(n_1753));

	AOI21X1 i_1837229(
		.A0(n_923),
		.A1(n_1753),
		.B0(n_1752),
		.Y(n_1754));

	NOR2BX1 i_847131(
		.AN(op_a[20]),
		.B(op_b[20]),
		.Y(n_1755));

	NOR2BX1 i_837130(
		.AN(op_a[19]),
		.B(op_b[19]),
		.Y(n_1756));

	AOI21X1 i_1817227(
		.A0(n_925),
		.A1(n_1756),
		.B0(n_1755),
		.Y(n_1757));

	AND2X1 i_2157259(
		.A(n_923),
		.B(n_1485),
		.Y(n_1758));

	NOR2BX1 i_827129(
		.AN(op_a[18]),
		.B(op_b[18]),
		.Y(n_1760));

	NOR2BX1 i_817128(
		.AN(op_a[17]),
		.B(op_b[17]),
		.Y(n_1761));

	AOI21X1 i_1797225(
		.A0(n_927),
		.A1(n_1761),
		.B0(n_1760),
		.Y(n_1762));

	NOR2BX1 i_807127(
		.AN(op_a[16]),
		.B(op_b[16]),
		.Y(n_1763));

	NOR2BX1 i_797126(
		.AN(op_a[15]),
		.B(op_b[15]),
		.Y(n_1764));

	AOI21X1 i_1777223(
		.A0(n_929),
		.A1(n_1764),
		.B0(n_1763),
		.Y(n_1765));

	NAND2X1 i_2117255(
		.A(n_927),
		.B(n_1383),
		.Y(n_1766));

	NOR2BX1 i_787125(
		.AN(n_7270),
		.B(op_b[14]),
		.Y(n_1768));

	NOR2BX1 i_777124(
		.AN(op_a[13]),
		.B(op_b[13]),
		.Y(n_1769));

	AOI21X1 i_1757221(
		.A0(n_931),
		.A1(n_1769),
		.B0(n_1768),
		.Y(n_1770));

	NOR2BX1 i_767123(
		.AN(op_a[12]),
		.B(op_b[12]),
		.Y(n_1771));

	NOR2BX1 i_757122(
		.AN(op_a[11]),
		.B(op_b[11]),
		.Y(n_1772));

	AOI21X1 i_1737219(
		.A0(n_933),
		.A1(n_1772),
		.B0(n_1771),
		.Y(n_1773));

	NAND2X1 i_2077251(
		.A(n_931),
		.B(n_1286),
		.Y(n_1774));

	NOR2BX1 i_747121(
		.AN(n_7290),
		.B(op_b[10]),
		.Y(n_1776));

	NOR2BX1 i_737120(
		.AN(op_a[9]),
		.B(op_b[9]),
		.Y(n_1777));

	AOI21X1 i_1717217(
		.A0(n_935),
		.A1(n_1777),
		.B0(n_1776),
		.Y(n_1778));

	NOR2BX1 i_727119(
		.AN(op_a[8]),
		.B(op_b[8]),
		.Y(n_1779));

	NOR2BX1 i_717118(
		.AN(op_a[7]),
		.B(op_b[7]),
		.Y(n_1780));

	AOI21X1 i_1697215(
		.A0(n_937),
		.A1(n_1780),
		.B0(n_1779),
		.Y(n_1781));

	NAND2X1 i_2037247(
		.A(n_935),
		.B(n_1186),
		.Y(n_1782));

	NOR2BX1 i_707117(
		.AN(op_a[6]),
		.B(op_b[6]),
		.Y(n_1784));

	NAND2BX1 i_697116(
		.AN(op_b[5]),
		.B(op_a[5]),
		.Y(n_1785));

	OAI21XL i_1677213(
		.A0(n_1785),
		.A1(n_940),
		.B0(n_3074),
		.Y(n_1786));

	NOR2BX1 i_687115(
		.AN(op_a[4]),
		.B(op_b[4]),
		.Y(n_1787));

	NOR2BX1 i_677114(
		.AN(n_7302),
		.B(op_b[3]),
		.Y(n_1788));

	AOI21X1 i_1657211(
		.A0(n_942),
		.A1(n_1788),
		.B0(n_1787),
		.Y(n_1789));

	NAND2BX1 i_1997243(
		.AN(n_940),
		.B(n_1090),
		.Y(n_1790));

	NOR2BX1 i_667113(
		.AN(op_a[2]),
		.B(op_b[2]),
		.Y(n_1792));

	NOR2BX1 i_657112(
		.AN(op_a[1]),
		.B(op_b[1]),
		.Y(n_1793));

	AOI21X1 i_1637209(
		.A0(n_1068),
		.A1(n_1793),
		.B0(n_1792),
		.Y(n_1794));

	NAND2BX1 i_1617207(
		.AN(op_a[0]),
		.B(op_b[0]),
		.Y(n_1795));

	NAND2X1 i_2267266(
		.A(n_857),
		.B(n_1794),
		.Y(n_1797));

	NAND2X1 i_1977241(
		.A(n_942),
		.B(n_1045),
		.Y(n_1798));

	NOR2X1 i_531(
		.A(n_1790),
		.B(n_1798),
		.Y(n_1799));

	NAND2X1 i_2017245(
		.A(n_937),
		.B(n_1135),
		.Y(n_1800));

	NAND2X1 i_2057249(
		.A(n_933),
		.B(n_1237),
		.Y(n_1802));

	NAND2X1 i_2097253(
		.A(n_929),
		.B(n_1332),
		.Y(n_1804));

	NAND2X1 i_2137257(
		.A(n_925),
		.B(n_1434),
		.Y(n_1806));

	NAND2X1 i_2177261(
		.A(n_921),
		.B(n_1532),
		.Y(n_1808));

	NOR2X1 i_15(
		.A(n_1750),
		.B(n_1808),
		.Y(n_1809));

	AOI21X1 i_443(
		.A0(n_955),
		.A1(n_954),
		.B0(n_952),
		.Y(n_1810));

	NAND2X1 i_611415(
		.A(op_a[29]),
		.B(op_b[29]),
		.Y(n_1812));

	NAND2X1 i_601414(
		.A(op_a[28]),
		.B(op_b[28]),
		.Y(n_1813));

	NAND2X1 i_591413(
		.A(op_a[27]),
		.B(op_b[27]),
		.Y(n_1814));

	OAI21XL i_1561510(
		.A0(n_1814),
		.A1(n_1697),
		.B0(n_1813),
		.Y(n_1815));

	NOR2X1 i_12(
		.A(n_1650),
		.B(n_1697),
		.Y(n_1816));

	NAND2X1 i_581412(
		.A(op_a[26]),
		.B(op_b[26]),
		.Y(n_1817));

	NAND2X1 i_571411(
		.A(op_a[25]),
		.B(op_b[25]),
		.Y(n_1818));

	OAI21XL i_1541508(
		.A0(n_1700),
		.A1(n_1818),
		.B0(n_1817),
		.Y(n_1819));

	NAND2X1 i_561410(
		.A(op_a[24]),
		.B(op_b[24]),
		.Y(n_1820));

	NAND2X1 i_551409(
		.A(op_a[23]),
		.B(op_b[23]),
		.Y(n_1821));

	OAI21XL i_1521506(
		.A0(n_1544),
		.A1(n_1821),
		.B0(n_1820),
		.Y(n_1822));

	NOR2X1 i_185(
		.A(n_1700),
		.B(n_1592),
		.Y(n_1823));

	NAND2X1 i_541408(
		.A(op_a[22]),
		.B(op_b[22]),
		.Y(n_1825));

	NAND2X1 i_531407(
		.A(op_a[21]),
		.B(op_b[21]),
		.Y(n_1826));

	OAI21XL i_1501504(
		.A0(n_1497),
		.A1(n_1826),
		.B0(n_1825),
		.Y(n_1827));

	NAND2X1 i_521406(
		.A(op_a[20]),
		.B(op_b[20]),
		.Y(n_1828));

	NAND2X1 i_511405(
		.A(op_a[19]),
		.B(op_b[19]),
		.Y(n_1829));

	OAI21XL i_1481502(
		.A0(n_1446),
		.A1(n_1829),
		.B0(n_1828),
		.Y(n_1830));

	NOR2X1 i_181(
		.A(n_1497),
		.B(n_1492),
		.Y(n_1831));

	NAND2X1 i_501404(
		.A(op_a[18]),
		.B(op_b[18]),
		.Y(n_1833));

	NAND2X1 i_491403(
		.A(op_a[17]),
		.B(op_b[17]),
		.Y(n_1834));

	OAI21XL i_1461500(
		.A0(n_1395),
		.A1(n_1834),
		.B0(n_1833),
		.Y(n_1835));

	NAND2X1 i_481402(
		.A(op_a[16]),
		.B(op_b[16]),
		.Y(n_1836));

	NAND2X1 i_471401(
		.A(op_a[15]),
		.B(op_b[15]),
		.Y(n_1837));

	OAI21XL i_1441498(
		.A0(n_1344),
		.A1(n_1837),
		.B0(n_1836),
		.Y(n_1838));

	NOR2X1 i_177(
		.A(n_1395),
		.B(n_1390),
		.Y(n_1839));

	NAND2X1 i_461400(
		.A(n_7270),
		.B(op_b[14]),
		.Y(n_1841));

	NAND2X1 i_451399(
		.A(op_a[13]),
		.B(op_b[13]),
		.Y(n_1842));

	OAI21XL i_1421496(
		.A0(n_1297),
		.A1(n_1842),
		.B0(n_1841),
		.Y(n_1843));

	NAND2X1 i_441398(
		.A(op_a[12]),
		.B(op_b[12]),
		.Y(n_1844));

	NAND2X1 i_431397(
		.A(op_a[11]),
		.B(op_b[11]),
		.Y(n_1845));

	OAI21XL i_1401494(
		.A0(n_1249),
		.A1(n_1845),
		.B0(n_1844),
		.Y(n_1846));

	NOR2X1 i_173(
		.A(n_1297),
		.B(n_1293),
		.Y(n_1847));

	NAND2X1 i_421396(
		.A(n_7290),
		.B(op_b[10]),
		.Y(n_1849));

	NAND2X1 i_411395(
		.A(op_a[9]),
		.B(op_b[9]),
		.Y(n_1850));

	OAI21XL i_1381492(
		.A0(n_1198),
		.A1(n_1850),
		.B0(n_1849),
		.Y(n_1851));

	NAND2X1 i_401394(
		.A(op_a[8]),
		.B(op_b[8]),
		.Y(n_1852));

	NAND2X1 i_391393(
		.A(op_a[7]),
		.B(op_b[7]),
		.Y(n_1853));

	OAI21XL i_1361490(
		.A0(n_1147),
		.A1(n_1853),
		.B0(n_1852),
		.Y(n_1854));

	NOR2X1 i_169(
		.A(n_1198),
		.B(n_1193),
		.Y(n_1855));

	NAND2X1 i_381392(
		.A(op_a[6]),
		.B(op_b[6]),
		.Y(n_1857));

	NAND2X1 i_371391(
		.A(op_a[5]),
		.B(op_b[5]),
		.Y(n_1858));

	OAI21XL i_1341488(
		.A0(n_1100),
		.A1(n_1858),
		.B0(n_1857),
		.Y(n_1859));

	NAND2X1 i_361390(
		.A(op_a[4]),
		.B(op_b[4]),
		.Y(n_1860));

	NAND2X1 i_351389(
		.A(n_7302),
		.B(op_b[3]),
		.Y(n_1861));

	OAI21XL i_1321486(
		.A0(n_1053),
		.A1(n_1861),
		.B0(n_1860),
		.Y(n_1862));

	NOR2X1 i_1651517(
		.A(n_1100),
		.B(n_1095),
		.Y(n_1863));

	NAND2X1 i_341388(
		.A(op_a[2]),
		.B(op_b[2]),
		.Y(n_1865));

	NAND2X1 i_331387(
		.A(op_a[1]),
		.B(op_b[1]),
		.Y(n_1866));

	OAI21XL i_1301484(
		.A0(n_1096),
		.A1(n_1866),
		.B0(n_1865),
		.Y(n_1867));

	NAND2X1 i_321386(
		.A(op_a[0]),
		.B(op_b[0]),
		.Y(n_1868));

	NOR2X1 i_498(
		.A(n_1096),
		.B(n_1072),
		.Y(n_1869));

	AOI21X1 i_192(
		.A0(n_1869),
		.A1(n_3085),
		.B0(n_1867),
		.Y(n_1870));

	NOR2X1 i_1631515(
		.A(n_1053),
		.B(n_1097),
		.Y(n_1871));

	NOR2X1 i_1671519(
		.A(n_1147),
		.B(n_1144),
		.Y(n_1873));

	NOR2X1 i_171(
		.A(n_1249),
		.B(n_1244),
		.Y(n_1875));

	NOR2X1 i_175(
		.A(n_1344),
		.B(n_1339),
		.Y(n_1877));

	NOR2X1 i_179(
		.A(n_1446),
		.B(n_1441),
		.Y(n_1879));

	NAND2X1 i_509(
		.A(n_1831),
		.B(n_1879),
		.Y(n_1880));

	NOR2X1 i_183(
		.A(n_1544),
		.B(n_1539),
		.Y(n_1881));

	NAND2X1 i_16(
		.A(n_1823),
		.B(n_1881),
		.Y(n_1882));

	OAI2BB1X1 i_406(
		.A0N(op_a[30]),
		.A1N(op_b[30]),
		.B0(n_915),
		.Y(n_1883));

	NOR2X1 i_11787(
		.A(op_a[0]),
		.B(op_a[1]),
		.Y(n_1885));

	NOR3X1 i_341819(
		.A(op_a[0]),
		.B(op_a[1]),
		.C(op_a[2]),
		.Y(n_1886));

	NOR2X1 i_26(
		.A(op_a[6]),
		.B(op_a[7]),
		.Y(n_1887));

	NOR2X1 i_25(
		.A(op_a[4]),
		.B(op_a[5]),
		.Y(n_1888));

	NAND4BXL i_711854(
		.AN(n_7302),
		.B(n_1888),
		.C(n_1887),
		.D(n_1886),
		.Y(n_1891));

	NOR2X1 i_27(
		.A(op_a[8]),
		.B(op_a[9]),
		.Y(n_1892));

	NOR2X1 i_28(
		.A(n_7290),
		.B(op_a[11]),
		.Y(n_1893));

	NAND3BX1 i_1071887(
		.AN(n_1891),
		.B(n_1892),
		.C(n_1893),
		.Y(n_1895));

	NOR2X1 i_30(
		.A(op_a[13]),
		.B(n_7270),
		.Y(n_1896));

	NOR4BX1 i_1111891(
		.AN(n_1896),
		.B(op_a[12]),
		.C(op_a[15]),
		.D(n_1895),
		.Y(n_1899));

	NOR2X1 i_24(
		.A(op_a[16]),
		.B(op_a[17]),
		.Y(n_1900));

	NOR2X1 i_31(
		.A(op_a[18]),
		.B(op_a[19]),
		.Y(n_1901));

	NAND3X1 i_1471921(
		.A(n_1900),
		.B(n_1901),
		.C(n_1899),
		.Y(n_1903));

	NOR2X1 i_29(
		.A(op_a[22]),
		.B(op_a[23]),
		.Y(n_1904));

	NOR2X1 i_32(
		.A(op_a[20]),
		.B(op_a[21]),
		.Y(n_1905));

	NOR4BX1 i_1511925(
		.AN(n_1904),
		.B(op_a[20]),
		.C(op_a[21]),
		.D(n_1903),
		.Y(n_1907));

	NOR2X1 i_20(
		.A(op_a[26]),
		.B(op_a[27]),
		.Y(n_1908));

	NOR2X1 i_21(
		.A(op_a[24]),
		.B(op_a[25]),
		.Y(n_1909));

	NAND3X1 i_1551929(
		.A(n_1909),
		.B(n_1908),
		.C(n_1907),
		.Y(n_1911));

	NOR2X1 i_22(
		.A(op_a[28]),
		.B(op_a[29]),
		.Y(n_1912));

	NAND2X1 i_8(
		.A(ovm),
		.B(n_166),
		.Y(n_1915));

	NAND3X1 i_1095(
		.A(cmd[0]),
		.B(cmd[2]),
		.C(n_1736),
		.Y(n_1917));

	NOR2BX1 i_3(
		.AN(op_a[31]),
		.B(n_1917),
		.Y(n_1918));

	NOR2X1 i_459(
		.A(n_7302),
		.B(op_a[6]),
		.Y(n_1919));

	NAND3X1 i_701853(
		.A(n_1919),
		.B(n_1888),
		.C(n_1886),
		.Y(n_1921));

	NOR4BX1 i_1061886(
		.AN(n_1892),
		.B(op_a[7]),
		.C(n_7290),
		.D(n_1921),
		.Y(n_1924));

	NOR4X1 i_464(
		.A(op_a[11]),
		.B(op_a[12]),
		.C(op_a[13]),
		.D(n_7270),
		.Y(n_1926));

	NAND2X1 i_1101890(
		.A(n_1926),
		.B(n_1924),
		.Y(n_1927));

	NOR4BX1 i_1461920(
		.AN(n_1900),
		.B(op_a[15]),
		.C(op_a[18]),
		.D(n_1927),
		.Y(n_1930));

	NOR4X1 i_468(
		.A(op_a[19]),
		.B(op_a[22]),
		.C(op_a[20]),
		.D(op_a[21]),
		.Y(n_1932));

	NAND2X1 i_1501924(
		.A(n_1932),
		.B(n_1930),
		.Y(n_1933));

	NOR4BX1 i_1541928(
		.AN(n_1909),
		.B(op_a[23]),
		.C(op_a[26]),
		.D(n_1933),
		.Y(n_1936));

	NOR4X1 i_561(
		.A(op_a[27]),
		.B(op_a[30]),
		.C(op_a[28]),
		.D(op_a[29]),
		.Y(n_1938));

	NAND3BX1 i_1088(
		.AN(cmd[2]),
		.B(cmd[1]),
		.C(cmd[0]),
		.Y(n_1942));

	NAND3BX1 i_1098(
		.AN(cmd[0]),
		.B(cmd[2]),
		.C(cmd[1]),
		.Y(n_1944));

	AND2X1 i_1100(
		.A(cmd[0]),
		.B(cmd[1]),
		.Y(n_1946));

	AOI22X1 i_564(
		.A0(op_b[31]),
		.A1(n_1946),
		.B0(n_963),
		.B1(op_a[31]),
		.Y(n_1947));

	OAI211X1 i_566(
		.A0(n_964),
		.A1(n_1740),
		.B0(n_967),
		.C0(n_1947),
		.Y(n_1949));

	AOI21X1 i_11(
		.A0(op_b[31]),
		.A1(n_3095),
		.B0(n_970),
		.Y(n_1950));

	NAND4BXL i_578(
		.AN(n_974),
		.B(n_1944),
		.C(n_1917),
		.D(n_7356),
		.Y(n_1955));

	AOI221X1 i_586(
		.A0(n_978),
		.A1(op_b[0]),
		.B0(n_7320),
		.B1(n_3085),
		.C0(n_6909),
		.Y(n_1957));

	NAND2X1 i_39(
		.A(n_3075),
		.B(n_3065),
		.Y(n_1959));

	NAND2X1 i_42(
		.A(op_a[31]),
		.B(op_a[0]),
		.Y(n_1961));

	AOI21X1 i_593(
		.A0(n_1961),
		.A1(op_a[1]),
		.B0(n_986),
		.Y(n_1962));

	AOI222X1 i_607(
		.A0(n_7320),
		.A1(n_3083),
		.B0(op_a[1]),
		.B1(n_3063),
		.C0(n_1946),
		.C1(op_b[1]),
		.Y(n_1965));

	OAI21XL i_608(
		.A0(n_1072),
		.A1(n_1942),
		.B0(n_1965),
		.Y(n_1966));

	AOI211X1 i_610(
		.A0(n_993),
		.A1(n_7341),
		.B0(n_1966),
		.C0(n_999),
		.Y(n_1968));

	OAI31X1 i_611(
		.A0(n_1959),
		.A1(n_1795),
		.A2(n_6939),
		.B0(n_1968),
		.Y(n_1969));

	NAND2BX1 i_45(
		.AN(n_1792),
		.B(n_1068),
		.Y(n_1970));

	OAI21XL i_1627208(
		.A0(op_b[0]),
		.A1(n_1136),
		.B0(n_3075),
		.Y(n_1971));

	NAND2BX1 i_2257265(
		.AN(n_1971),
		.B(n_856),
		.Y(n_1972));

	OAI21XL i_48(
		.A0(op_a[0]),
		.A1(op_a[1]),
		.B0(op_a[31]),
		.Y(n_1974));

	AOI21X1 i_618(
		.A0(n_1974),
		.A1(op_a[2]),
		.B0(n_1006),
		.Y(n_1975));

	OAI21XL i_1291483(
		.A0(n_1072),
		.A1(n_1868),
		.B0(n_1866),
		.Y(n_1976));

	NOR2X1 i_47(
		.A(n_1096),
		.B(n_3084),
		.Y(n_1977));

	AOI222X1 i_633(
		.A0(n_7320),
		.A1(n_3084),
		.B0(op_a[2]),
		.B1(n_3063),
		.C0(n_1946),
		.C1(op_b[2]),
		.Y(n_1979));

	OAI21XL i_634(
		.A0(n_1096),
		.A1(n_1942),
		.B0(n_1979),
		.Y(n_1980));

	AOI211X1 i_636(
		.A0(n_1014),
		.A1(n_7341),
		.B0(n_1980),
		.C0(n_1020),
		.Y(n_1982));

	OAI31X1 i_637(
		.A0(n_1970),
		.A1(n_7387),
		.A2(n_1972),
		.B0(n_1982),
		.Y(n_1983));

	NAND2BX1 i_51(
		.AN(n_1788),
		.B(n_1045),
		.Y(n_1984));

	NAND2X1 i_54(
		.A(op_a[31]),
		.B(n_3067),
		.Y(n_1986));

	AOI21X1 i_643(
		.A0(n_7302),
		.A1(n_1986),
		.B0(n_1026),
		.Y(n_1987));

	NOR2X1 i_53(
		.A(n_1097),
		.B(n_3081),
		.Y(n_1988));

	AOI222X1 i_657(
		.A0(n_7320),
		.A1(n_3081),
		.B0(n_7302),
		.B1(n_3063),
		.C0(n_1946),
		.C1(op_b[3]),
		.Y(n_1990));

	OAI21XL i_658(
		.A0(n_1097),
		.A1(n_7356),
		.B0(n_1990),
		.Y(n_1991));

	AOI211X1 i_660(
		.A0(n_1033),
		.A1(n_7341),
		.B0(n_1991),
		.C0(n_1039),
		.Y(n_1993));

	OAI31X1 i_661(
		.A0(n_1984),
		.A1(n_1797),
		.A2(n_6939),
		.B0(n_1993),
		.Y(n_1994));

	NAND2BX1 i_57(
		.AN(n_1787),
		.B(n_942),
		.Y(n_1995));

	AOI21X1 i_1647210(
		.A0(n_1045),
		.A1(n_1792),
		.B0(n_1788),
		.Y(n_1996));

	NAND2X1 i_1967240(
		.A(n_1045),
		.B(n_1068),
		.Y(n_1997));

	AOI31X1 i_2277267(
		.A0(n_1971),
		.A1(n_1045),
		.A2(n_1068),
		.B0(n_3087),
		.Y(n_1998));

	OAI21XL i_17(
		.A0(n_7302),
		.A1(n_3067),
		.B0(op_a[31]),
		.Y(n_2000));

	AOI21X1 i_671(
		.A0(n_2000),
		.A1(op_a[4]),
		.B0(n_1048),
		.Y(n_2001));

	OAI21XL i_1311485(
		.A0(n_1097),
		.A1(n_1865),
		.B0(n_1861),
		.Y(n_2002));

	NOR2X1 i_674(
		.A(n_1097),
		.B(n_1096),
		.Y(n_2003));

	AOI21X1 i_193(
		.A0(n_1976),
		.A1(n_2003),
		.B0(n_2002),
		.Y(n_2004));

	NOR2X1 i_59(
		.A(n_1053),
		.B(n_3082),
		.Y(n_2005));

	AOI222X1 i_687(
		.A0(n_7320),
		.A1(n_3082),
		.B0(op_a[4]),
		.B1(n_3063),
		.C0(n_1946),
		.C1(op_b[4]),
		.Y(n_2007));

	OAI21XL i_688(
		.A0(n_1053),
		.A1(n_7356),
		.B0(n_2007),
		.Y(n_2008));

	AOI211X1 i_690(
		.A0(n_1057),
		.A1(n_7341),
		.B0(n_2008),
		.C0(n_1063),
		.Y(n_2010));

	OAI31X1 i_691(
		.A0(n_1137),
		.A1(n_1995),
		.A2(n_6939),
		.B0(n_2010),
		.Y(n_2011));

	OAI21XL i_2287268(
		.A0(n_1798),
		.A1(n_1794),
		.B0(n_1789),
		.Y(n_2013));

	NOR2X1 i_699(
		.A(op_a[2]),
		.B(n_7302),
		.Y(n_2016));

	NOR4BX1 i_681851(
		.AN(n_1885),
		.B(op_a[2]),
		.C(n_7302),
		.D(op_a[4]),
		.Y(n_2017));

	NAND2BX1 i_65(
		.AN(n_2017),
		.B(op_a[31]),
		.Y(n_2018));

	AOI21X1 i_702(
		.A0(op_a[5]),
		.A1(n_2018),
		.B0(n_1070),
		.Y(n_2019));

	AOI21X1 i_194(
		.A0(n_1867),
		.A1(n_1871),
		.B0(n_1862),
		.Y(n_2020));

	NOR2X1 i_64(
		.A(n_1095),
		.B(n_3079),
		.Y(n_2021));

	AOI222X1 i_718(
		.A0(n_7320),
		.A1(n_3079),
		.B0(op_a[5]),
		.B1(n_3063),
		.C0(n_1946),
		.C1(op_b[5]),
		.Y(n_2023));

	OAI221XL i_720(
		.A0(n_1095),
		.A1(n_7356),
		.B0(n_1078),
		.B1(n_3095),
		.C0(n_2023),
		.Y(n_2025));

	NAND2BX1 i_68(
		.AN(n_940),
		.B(n_3074),
		.Y(n_2028));

	NAND2X1 i_1667212(
		.A(n_1089),
		.B(n_1785),
		.Y(n_2029));

	NAND3X1 i_691852(
		.A(n_1888),
		.B(n_2016),
		.C(n_1885),
		.Y(n_2035));

	NAND2X1 i_72(
		.A(n_2035),
		.B(op_a[31]),
		.Y(n_2036));

	AOI21X1 i_733(
		.A0(n_2036),
		.A1(op_a[6]),
		.B0(n_1092),
		.Y(n_2037));

	OAI21XL i_1331487(
		.A0(n_1095),
		.A1(n_1860),
		.B0(n_1858),
		.Y(n_2038));

	NOR2X1 i_1641516(
		.A(n_1095),
		.B(n_1053),
		.Y(n_2039));

	AOI21X1 i_195(
		.A0(n_2002),
		.A1(n_2039),
		.B0(n_2038),
		.Y(n_2040));

	NOR2X1 i_70(
		.A(n_1100),
		.B(n_3080),
		.Y(n_2042));

	AOI222X1 i_750(
		.A0(n_7320),
		.A1(n_3080),
		.B0(op_a[6]),
		.B1(n_3063),
		.C0(n_1946),
		.C1(op_b[6]),
		.Y(n_2044));

	OAI21XL i_751(
		.A0(n_1100),
		.A1(n_1942),
		.B0(n_2044),
		.Y(n_2045));

	AOI211X1 i_753(
		.A0(n_1104),
		.A1(n_7341),
		.B0(n_2045),
		.C0(n_1110),
		.Y(n_2047));

	OAI31X1 i_754(
		.A0(n_2028),
		.A1(n_7387),
		.A2(n_1187),
		.B0(n_2047),
		.Y(n_2048));

	NAND2BX1 i_75(
		.AN(n_1780),
		.B(n_1135),
		.Y(n_2049));

	NAND2X1 i_78(
		.A(n_1921),
		.B(op_a[31]),
		.Y(n_2051));

	AOI21X1 i_760(
		.A0(n_2051),
		.A1(op_a[7]),
		.B0(n_1116),
		.Y(n_2052));

	NOR2X1 i_77(
		.A(n_1144),
		.B(n_3078),
		.Y(n_2053));

	AOI222X1 i_774(
		.A0(n_7320),
		.A1(n_3078),
		.B0(op_a[7]),
		.B1(n_3063),
		.C0(n_1946),
		.C1(op_b[7]),
		.Y(n_2055));

	OAI21XL i_775(
		.A0(n_1144),
		.A1(n_7356),
		.B0(n_2055),
		.Y(n_2056));

	AOI211X1 i_777(
		.A0(n_1123),
		.A1(n_7341),
		.B0(n_2056),
		.C0(n_1129),
		.Y(n_2058));

	OAI31X1 i_778(
		.A0(n_2049),
		.A1(n_7387),
		.A2(n_3076),
		.B0(n_2058),
		.Y(n_2059));

	NAND2BX1 i_82(
		.AN(n_1779),
		.B(n_937),
		.Y(n_2060));

	AOI21X1 i_1687214(
		.A0(n_1135),
		.A1(n_1784),
		.B0(n_1780),
		.Y(n_2061));

	NOR2BX1 i_2007244(
		.AN(n_1135),
		.B(n_940),
		.Y(n_2062));

	OAI21XL i_1351489(
		.A0(n_1144),
		.A1(n_1857),
		.B0(n_1853),
		.Y(n_2066));

	NOR2X1 i_1661518(
		.A(n_1144),
		.B(n_1100),
		.Y(n_2067));

	AOI21X1 i_83(
		.A0(op_a[8]),
		.A1(op_b[8]),
		.B0(n_1147),
		.Y(n_2070));

	OAI21XL i_0(
		.A0(op_a[31]),
		.A1(n_1917),
		.B0(n_1944),
		.Y(n_2071));

	OAI211X1 i_804(
		.A0(op_a[8]),
		.A1(n_7313),
		.B0(op_b[8]),
		.C0(n_7317),
		.Y(n_2072));

	OAI221XL i_806(
		.A0(n_1147),
		.A1(n_1942),
		.B0(n_1150),
		.B1(n_3068),
		.C0(n_2072),
		.Y(n_2074));

	AOI221X1 i_808(
		.A0(n_7338),
		.A1(op_a[8]),
		.B0(n_1151),
		.B1(n_7341),
		.C0(n_2074),
		.Y(n_2076));

	OAI31X1 i_809(
		.A0(n_2060),
		.A1(n_6939),
		.A2(n_1238),
		.B0(n_2076),
		.Y(n_2077));

	NAND2BX1 i_87(
		.AN(n_1777),
		.B(n_1186),
		.Y(n_2079));

	AOI31X1 i_2327272(
		.A0(n_937),
		.A1(n_1786),
		.A2(n_1135),
		.B0(n_3073),
		.Y(n_2080));

	AOI21X1 i_198(
		.A0(n_1859),
		.A1(n_1873),
		.B0(n_1854),
		.Y(n_2083));

	AOI21X1 i_88(
		.A0(op_a[9]),
		.A1(op_b[9]),
		.B0(n_1193),
		.Y(n_2085));

	NOR4X1 i_818(
		.A(op_a[6]),
		.B(op_a[7]),
		.C(op_a[5]),
		.D(op_a[8]),
		.Y(n_2087));

	NAND2X1 i_1041884(
		.A(n_2087),
		.B(n_2017),
		.Y(n_2088));

	OAI211X1 i_834(
		.A0(op_a[9]),
		.A1(n_7313),
		.B0(op_b[9]),
		.C0(cmd[1]),
		.Y(n_2089));

	OAI221XL i_836(
		.A0(n_1193),
		.A1(n_1942),
		.B0(n_1173),
		.B1(n_3068),
		.C0(n_2089),
		.Y(n_2091));

	AOI221X1 i_838(
		.A0(n_7338),
		.A1(op_a[9]),
		.B0(n_1174),
		.B1(n_7341),
		.C0(n_2091),
		.Y(n_2093));

	OAI31X1 i_839(
		.A0(n_2079),
		.A1(n_6939),
		.A2(n_1264),
		.B0(n_2093),
		.Y(n_2094));

	NAND2BX1 i_92(
		.AN(n_1776),
		.B(n_935),
		.Y(n_2096));

	AOI21X1 i_1707216(
		.A0(n_1186),
		.A1(n_1779),
		.B0(n_1777),
		.Y(n_2097));

	NAND2X1 i_2027246(
		.A(n_1186),
		.B(n_937),
		.Y(n_2098));

	OAI21XL i_1371491(
		.A0(n_1193),
		.A1(n_1852),
		.B0(n_1850),
		.Y(n_2102));

	NOR2X1 i_168(
		.A(n_1193),
		.B(n_1147),
		.Y(n_2103));

	AOI21X1 i_93(
		.A0(n_7290),
		.A1(op_b[10]),
		.B0(n_1198),
		.Y(n_2106));

	NOR4BX1 i_1051885(
		.AN(n_1887),
		.B(op_a[8]),
		.C(op_a[9]),
		.D(n_2035),
		.Y(n_2108));

	OAI211X1 i_866(
		.A0(n_7290),
		.A1(n_7313),
		.B0(op_b[10]),
		.C0(n_7320),
		.Y(n_2109));

	OAI221XL i_868(
		.A0(n_1198),
		.A1(n_1942),
		.B0(n_1201),
		.B1(n_6911),
		.C0(n_2109),
		.Y(n_2111));

	AOI221X1 i_870(
		.A0(n_7338),
		.A1(n_7290),
		.B0(n_1202),
		.B1(n_7341),
		.C0(n_2111),
		.Y(n_2113));

	OAI31X1 i_871(
		.A0(n_2096),
		.A1(n_6939),
		.A2(n_1287),
		.B0(n_2113),
		.Y(n_2114));

	NAND2BX1 i_97(
		.AN(n_1772),
		.B(n_1237),
		.Y(n_2116));

	AOI21X1 i_98(
		.A0(op_a[11]),
		.A1(op_b[11]),
		.B0(n_1244),
		.Y(n_2118));

	OAI211X1 i_896(
		.A0(op_a[11]),
		.A1(n_7313),
		.B0(op_b[11]),
		.C0(n_7317),
		.Y(n_2119));

	OAI221XL i_898(
		.A0(n_1244),
		.A1(n_1942),
		.B0(n_1224),
		.B1(n_3068),
		.C0(n_2119),
		.Y(n_2121));

	AOI221X1 i_900(
		.A0(n_7338),
		.A1(op_a[11]),
		.B0(n_1225),
		.B1(n_6904),
		.C0(n_2121),
		.Y(n_2123));

	OAI31X1 i_901(
		.A0(n_2116),
		.A1(n_6939),
		.A2(n_943),
		.B0(n_2123),
		.Y(n_2124));

	NAND2BX1 i_102(
		.AN(n_1771),
		.B(n_933),
		.Y(n_2126));

	AOI21X1 i_1727218(
		.A0(n_1237),
		.A1(n_1776),
		.B0(n_1772),
		.Y(n_2127));

	NAND2X1 i_2047248(
		.A(n_1237),
		.B(n_935),
		.Y(n_2128));

	OAI21XL i_1391493(
		.A0(n_1244),
		.A1(n_1849),
		.B0(n_1845),
		.Y(n_2132));

	NOR2X1 i_170(
		.A(n_1244),
		.B(n_1198),
		.Y(n_2133));

	AOI21X1 i_104(
		.A0(op_a[12]),
		.A1(op_b[12]),
		.B0(n_1249),
		.Y(n_2136));

	OAI211X1 i_928(
		.A0(op_a[12]),
		.A1(n_7313),
		.B0(op_b[12]),
		.C0(n_7317),
		.Y(n_2137));

	OAI221XL i_930(
		.A0(n_1249),
		.A1(n_1942),
		.B0(n_1252),
		.B1(n_3068),
		.C0(n_2137),
		.Y(n_2139));

	AOI221X1 i_932(
		.A0(n_7338),
		.A1(op_a[12]),
		.B0(n_1253),
		.B1(n_7341),
		.C0(n_2139),
		.Y(n_2141));

	OAI31X1 i_933(
		.A0(n_2126),
		.A1(n_6939),
		.A2(n_1334),
		.B0(n_2141),
		.Y(n_2142));

	NAND2BX1 i_108(
		.AN(n_1769),
		.B(n_1286),
		.Y(n_2144));

	AOI21X1 i_109(
		.A0(op_a[13]),
		.A1(op_b[13]),
		.B0(n_1293),
		.Y(n_2150));

	NOR4BX1 i_1081888(
		.AN(n_1893),
		.B(op_a[9]),
		.C(op_a[12]),
		.D(n_2088),
		.Y(n_2153));

	OAI211X1 i_960(
		.A0(op_a[13]),
		.A1(n_7313),
		.B0(op_b[13]),
		.C0(n_7317),
		.Y(n_2154));

	OAI221XL i_962(
		.A0(n_1293),
		.A1(n_6901),
		.B0(n_1273),
		.B1(n_3068),
		.C0(n_2154),
		.Y(n_2156));

	AOI221X1 i_964(
		.A0(n_6906),
		.A1(op_a[13]),
		.B0(n_1274),
		.B1(n_7341),
		.C0(n_2156),
		.Y(n_2158));

	OAI31X1 i_965(
		.A0(n_2144),
		.A1(n_6939),
		.A2(n_1360),
		.B0(n_2158),
		.Y(n_2159));

	NAND2BX1 i_113(
		.AN(n_1768),
		.B(n_931),
		.Y(n_2161));

	AOI21X1 i_1747220(
		.A0(n_1286),
		.A1(n_1771),
		.B0(n_1769),
		.Y(n_2162));

	NAND2X1 i_2067250(
		.A(n_1286),
		.B(n_933),
		.Y(n_2163));

	OAI21XL i_1411495(
		.A0(n_1293),
		.A1(n_1844),
		.B0(n_1842),
		.Y(n_2167));

	NOR2X1 i_172(
		.A(n_1293),
		.B(n_1249),
		.Y(n_2168));

	AOI21X1 i_114(
		.A0(n_7270),
		.A1(op_b[14]),
		.B0(n_1297),
		.Y(n_2171));

	NOR4BBX1 i_1091889(
		.AN(n_1893),
		.BN(n_2108),
		.C(op_a[12]),
		.D(op_a[13]),
		.Y(n_2174));

	OAI211X1 i_994(
		.A0(n_7270),
		.A1(n_7313),
		.B0(op_b[14]),
		.C0(n_7320),
		.Y(n_2175));

	OAI221XL i_996(
		.A0(n_1297),
		.A1(n_6901),
		.B0(n_1300),
		.B1(n_3068),
		.C0(n_2175),
		.Y(n_2177));

	AOI221X1 i_998(
		.A0(n_6906),
		.A1(n_7270),
		.B0(n_1301),
		.B1(n_7341),
		.C0(n_2177),
		.Y(n_2179));

	OAI31X1 i_999(
		.A0(n_2161),
		.A1(n_6939),
		.A2(n_1385),
		.B0(n_2179),
		.Y(n_2180));

	NAND2BX1 i_118(
		.AN(n_1764),
		.B(n_1332),
		.Y(n_2182));

	AOI21X1 i_119(
		.A0(op_a[15]),
		.A1(op_b[15]),
		.B0(n_1339),
		.Y(n_2184));

	OAI211X1 i_1018(
		.A0(op_a[15]),
		.A1(n_7313),
		.B0(op_b[15]),
		.C0(n_7317),
		.Y(n_2185));

	OAI221XL i_1020(
		.A0(n_1339),
		.A1(n_6901),
		.B0(n_1319),
		.B1(n_3068),
		.C0(n_2185),
		.Y(n_2187));

	AOI221X1 i_1022(
		.A0(n_7338),
		.A1(op_a[15]),
		.B0(n_1320),
		.B1(n_6904),
		.C0(n_2187),
		.Y(n_2189));

	OAI31X1 i_1023(
		.A0(n_2182),
		.A1(n_7323),
		.A2(n_1411),
		.B0(n_2189),
		.Y(n_2190));

	NAND2BX1 i_123(
		.AN(n_1763),
		.B(n_929),
		.Y(n_2192));

	AOI21X1 i_1767222(
		.A0(n_1332),
		.A1(n_1768),
		.B0(n_1764),
		.Y(n_2193));

	NAND2X1 i_2087252(
		.A(n_1332),
		.B(n_931),
		.Y(n_2194));

	OAI21XL i_1431497(
		.A0(n_1339),
		.A1(n_1841),
		.B0(n_1837),
		.Y(n_2198));

	NOR2X1 i_174(
		.A(n_1339),
		.B(n_1297),
		.Y(n_2199));

	AOI21X1 i_124(
		.A0(op_a[16]),
		.A1(op_b[16]),
		.B0(n_1344),
		.Y(n_2202));

	OAI211X1 i_1051(
		.A0(op_a[16]),
		.A1(n_7313),
		.B0(op_b[16]),
		.C0(n_7317),
		.Y(n_2203));

	OAI221XL i_1053(
		.A0(n_1344),
		.A1(n_6901),
		.B0(n_1347),
		.B1(n_6911),
		.C0(n_2203),
		.Y(n_2205));

	AOI221X1 i_1055(
		.A0(n_7338),
		.A1(op_a[16]),
		.B0(n_1348),
		.B1(n_6904),
		.C0(n_2205),
		.Y(n_2207));

	OAI31X1 i_1056(
		.A0(n_2192),
		.A1(n_7323),
		.A2(n_1436),
		.B0(n_2207),
		.Y(n_2208));

	NAND2BX1 i_128(
		.AN(n_1761),
		.B(n_1383),
		.Y(n_2210));

	AOI21X1 i_129(
		.A0(op_a[17]),
		.A1(op_b[17]),
		.B0(n_1390),
		.Y(n_2216));

	NOR4X1 i_1067(
		.A(op_a[13]),
		.B(n_7270),
		.C(op_a[15]),
		.D(op_a[16]),
		.Y(n_2218));

	NAND2X1 i_1441918(
		.A(n_2218),
		.B(n_2153),
		.Y(n_2219));

	OAI211X1 i_1089(
		.A0(op_a[17]),
		.A1(n_7313),
		.B0(op_b[17]),
		.C0(n_7317),
		.Y(n_2220));

	OAI221XL i_1091(
		.A0(n_1390),
		.A1(n_6901),
		.B0(n_1370),
		.B1(n_6911),
		.C0(n_2220),
		.Y(n_2222));

	AOI221X1 i_1094(
		.A0(n_7338),
		.A1(op_a[17]),
		.B0(n_1371),
		.B1(n_6904),
		.C0(n_2222),
		.Y(n_2224));

	OAI31X1 i_1096(
		.A0(n_2210),
		.A1(n_7323),
		.A2(n_1462),
		.B0(n_2224),
		.Y(n_2225));

	NAND2BX1 i_133(
		.AN(n_1760),
		.B(n_927),
		.Y(n_2227));

	AOI21X1 i_1787224(
		.A0(n_1383),
		.A1(n_1763),
		.B0(n_1761),
		.Y(n_2228));

	NAND2X1 i_2107254(
		.A(n_1383),
		.B(n_929),
		.Y(n_2229));

	OAI21XL i_1451499(
		.A0(n_1390),
		.A1(n_1836),
		.B0(n_1834),
		.Y(n_2233));

	NOR2X1 i_176(
		.A(n_1390),
		.B(n_1344),
		.Y(n_2234));

	AOI21X1 i_134(
		.A0(op_a[18]),
		.A1(op_b[18]),
		.B0(n_1395),
		.Y(n_2237));

	NOR4X1 i_1111(
		.A(op_a[16]),
		.B(op_a[17]),
		.C(n_7270),
		.D(op_a[15]),
		.Y(n_2239));

	OAI211X1 i_1132(
		.A0(op_a[18]),
		.A1(cmd[0]),
		.B0(op_b[18]),
		.C0(n_7320),
		.Y(n_2241));

	OAI221XL i_1134(
		.A0(n_1395),
		.A1(n_6901),
		.B0(n_1398),
		.B1(n_6911),
		.C0(n_2241),
		.Y(n_2243));

	AOI221X1 i_1137(
		.A0(n_7338),
		.A1(op_a[18]),
		.B0(n_1399),
		.B1(n_6904),
		.C0(n_2243),
		.Y(n_2245));

	OAI31X1 i_1138(
		.A0(n_2227),
		.A1(n_7323),
		.A2(n_1487),
		.B0(n_2245),
		.Y(n_2246));

	NAND2BX1 i_190(
		.AN(n_1756),
		.B(n_1434),
		.Y(n_2248));

	AOI21X1 i_191(
		.A0(op_a[19]),
		.A1(op_b[19]),
		.B0(n_1441),
		.Y(n_2250));

	OAI211X1 i_1168(
		.A0(op_a[19]),
		.A1(cmd[0]),
		.B0(op_b[19]),
		.C0(cmd[1]),
		.Y(n_2251));

	OAI221XL i_1170(
		.A0(n_1441),
		.A1(n_6901),
		.B0(n_1421),
		.B1(n_6911),
		.C0(n_2251),
		.Y(n_2253));

	AOI221X1 i_1173(
		.A0(n_6906),
		.A1(op_a[19]),
		.B0(n_1422),
		.B1(n_6904),
		.C0(n_2253),
		.Y(n_2255));

	OAI31X1 i_1174(
		.A0(n_2248),
		.A1(n_7323),
		.A2(n_946),
		.B0(n_2255),
		.Y(n_2256));

	NAND2BX1 i_222(
		.AN(n_1755),
		.B(n_925),
		.Y(n_2258));

	AOI21X1 i_1807226(
		.A0(n_1434),
		.A1(n_1760),
		.B0(n_1756),
		.Y(n_2259));

	NAND2X1 i_2127256(
		.A(n_1434),
		.B(n_927),
		.Y(n_2260));

	OAI21XL i_1471501(
		.A0(n_1441),
		.A1(n_1833),
		.B0(n_1829),
		.Y(n_2264));

	NOR2X1 i_178(
		.A(n_1441),
		.B(n_1395),
		.Y(n_2265));

	AOI21X1 i_224(
		.A0(op_a[20]),
		.A1(op_b[20]),
		.B0(n_1446),
		.Y(n_2268));

	OAI211X1 i_1206(
		.A0(op_a[20]),
		.A1(cmd[0]),
		.B0(op_b[20]),
		.C0(n_7317),
		.Y(n_2269));

	OAI221XL i_1209(
		.A0(n_1446),
		.A1(n_6901),
		.B0(n_1449),
		.B1(n_6911),
		.C0(n_2269),
		.Y(n_2271));

	AOI221X1 i_1211(
		.A0(n_6906),
		.A1(op_a[20]),
		.B0(n_1450),
		.B1(n_6904),
		.C0(n_2271),
		.Y(n_2273));

	OAI31X1 i_1212(
		.A0(n_2258),
		.A1(n_7323),
		.A2(n_1534),
		.B0(n_2273),
		.Y(n_2274));

	NAND2BX1 i_229(
		.AN(n_1753),
		.B(n_1485),
		.Y(n_2276));

	AOI21X1 i_230(
		.A0(op_a[21]),
		.A1(op_b[21]),
		.B0(n_1492),
		.Y(n_2282));

	NOR4BX1 i_1481922(
		.AN(n_1901),
		.B(op_a[17]),
		.C(op_a[20]),
		.D(n_2219),
		.Y(n_2285));

	OAI211X1 i_1245(
		.A0(op_a[21]),
		.A1(cmd[0]),
		.B0(op_b[21]),
		.C0(cmd[1]),
		.Y(n_2286));

	OAI221XL i_1247(
		.A0(n_1492),
		.A1(n_6901),
		.B0(n_1472),
		.B1(n_6911),
		.C0(n_2286),
		.Y(n_2288));

	AOI221X1 i_1249(
		.A0(n_6906),
		.A1(op_a[21]),
		.B0(n_1473),
		.B1(n_6904),
		.C0(n_2288),
		.Y(n_2290));

	OAI31X1 i_1250(
		.A0(n_2276),
		.A1(n_6939),
		.A2(n_1561),
		.B0(n_2290),
		.Y(n_2291));

	NAND2BX1 i_236(
		.AN(n_1752),
		.B(n_923),
		.Y(n_2293));

	AOI21X1 i_1827228(
		.A0(n_1485),
		.A1(n_1755),
		.B0(n_1753),
		.Y(n_2294));

	NAND2X1 i_2147258(
		.A(n_1485),
		.B(n_925),
		.Y(n_2295));

	OAI21XL i_1491503(
		.A0(n_1492),
		.A1(n_1828),
		.B0(n_1826),
		.Y(n_2299));

	NOR2X1 i_180(
		.A(n_1492),
		.B(n_1446),
		.Y(n_2300));

	AOI21X1 i_237(
		.A0(op_a[22]),
		.A1(op_b[22]),
		.B0(n_1497),
		.Y(n_2303));

	NAND4X1 i_1491923(
		.A(n_1905),
		.B(n_1901),
		.C(n_2239),
		.D(n_2174),
		.Y(n_2305));

	OAI211X1 i_1284(
		.A0(op_a[22]),
		.A1(cmd[0]),
		.B0(op_b[22]),
		.C0(cmd[1]),
		.Y(n_2306));

	OAI221XL i_1286(
		.A0(n_1497),
		.A1(n_6901),
		.B0(n_1500),
		.B1(n_6911),
		.C0(n_2306),
		.Y(n_2308));

	AOI221X1 i_1289(
		.A0(n_6906),
		.A1(op_a[22]),
		.B0(n_1501),
		.B1(n_6904),
		.C0(n_2308),
		.Y(n_2310));

	OAI31X1 i_1290(
		.A0(n_2293),
		.A1(n_6939),
		.A2(n_1587),
		.B0(n_2310),
		.Y(n_2311));

	NAND2BX1 i_242(
		.AN(n_1748),
		.B(n_1532),
		.Y(n_2313));

	AOI21X1 i_244(
		.A0(op_a[23]),
		.A1(op_b[23]),
		.B0(n_1539),
		.Y(n_2315));

	OAI211X1 i_1311(
		.A0(op_a[23]),
		.A1(cmd[0]),
		.B0(op_b[23]),
		.C0(cmd[1]),
		.Y(n_2316));

	OAI221XL i_1313(
		.A0(n_1539),
		.A1(n_6901),
		.B0(n_1519),
		.B1(n_6911),
		.C0(n_2316),
		.Y(n_2318));

	AOI221X1 i_1316(
		.A0(n_7338),
		.A1(op_a[23]),
		.B0(n_1520),
		.B1(n_6904),
		.C0(n_2318),
		.Y(n_2320));

	OAI31X1 i_1317(
		.A0(n_2313),
		.A1(n_7323),
		.A2(n_1612),
		.B0(n_2320),
		.Y(n_2321));

	NAND2BX1 i_249(
		.AN(n_1747),
		.B(n_921),
		.Y(n_2323));

	AOI21X1 i_1847230(
		.A0(n_1532),
		.A1(n_1752),
		.B0(n_1748),
		.Y(n_2324));

	NAND2X1 i_2167260(
		.A(n_1532),
		.B(n_923),
		.Y(n_2325));

	OAI21XL i_1511505(
		.A0(n_1539),
		.A1(n_1825),
		.B0(n_1821),
		.Y(n_2329));

	NOR2X1 i_182(
		.A(n_1539),
		.B(n_1497),
		.Y(n_2330));

	AOI21X1 i_250(
		.A0(op_a[24]),
		.A1(op_b[24]),
		.B0(n_1544),
		.Y(n_2333));

	OAI211X1 i_1349(
		.A0(op_a[24]),
		.A1(cmd[0]),
		.B0(op_b[24]),
		.C0(cmd[1]),
		.Y(n_2334));

	OAI221XL i_1352(
		.A0(n_1544),
		.A1(n_6901),
		.B0(n_1547),
		.B1(n_6911),
		.C0(n_2334),
		.Y(n_2336));

	AOI221X1 i_1354(
		.A0(n_7338),
		.A1(op_a[24]),
		.B0(n_1548),
		.B1(n_6904),
		.C0(n_2336),
		.Y(n_2338));

	OAI31X1 i_1355(
		.A0(n_2323),
		.A1(n_7323),
		.A2(n_1637),
		.B0(n_2338),
		.Y(n_2339));

	NAND2BX1 i_255(
		.AN(n_1745),
		.B(n_1585),
		.Y(n_2341));

	OAI21XL i_2487288(
		.A0(n_1754),
		.A1(n_1808),
		.B0(n_1749),
		.Y(n_2342));

	AOI31X1 i_4377415(
		.A0(n_1561),
		.A1(n_3071),
		.A2(n_1758),
		.B0(n_2342),
		.Y(n_2344));

	AOI21X1 i_214(
		.A0(n_1827),
		.A1(n_1881),
		.B0(n_1822),
		.Y(n_2346));

	AOI21X1 i_260(
		.A0(op_a[25]),
		.A1(op_b[25]),
		.B0(n_1592),
		.Y(n_2349));

	NOR4X1 i_1367(
		.A(op_a[22]),
		.B(op_a[23]),
		.C(op_a[21]),
		.D(op_a[24]),
		.Y(n_2351));

	NAND2X1 i_1521926(
		.A(n_2351),
		.B(n_2285),
		.Y(n_2352));

	OAI211X1 i_1399(
		.A0(op_a[25]),
		.A1(n_7313),
		.B0(op_b[25]),
		.C0(n_7320),
		.Y(n_2353));

	OAI221XL i_1401(
		.A0(n_1592),
		.A1(n_1942),
		.B0(n_1572),
		.B1(n_3068),
		.C0(n_2353),
		.Y(n_2355));

	AOI211X1 i_1403(
		.A0(n_7338),
		.A1(op_a[25]),
		.B0(n_2355),
		.C0(n_1579),
		.Y(n_2357));

	OAI31X1 i_1404(
		.A0(n_3093),
		.A1(n_2341),
		.A2(n_7323),
		.B0(n_2357),
		.Y(n_2358));

	NAND2BX1 i_264(
		.AN(n_1744),
		.B(n_1709),
		.Y(n_2360));

	AOI21X1 i_1867232(
		.A0(n_1585),
		.A1(n_1747),
		.B0(n_1745),
		.Y(n_2361));

	AND2X1 i_2187262(
		.A(n_1585),
		.B(n_921),
		.Y(n_2362));

	OAI21XL i_1531507(
		.A0(n_1592),
		.A1(n_1820),
		.B0(n_1818),
		.Y(n_2366));

	NOR2X1 i_184(
		.A(n_1592),
		.B(n_1544),
		.Y(n_2367));

	AOI21X1 i_265(
		.A0(op_a[26]),
		.A1(op_b[26]),
		.B0(n_1700),
		.Y(n_2370));

	NOR4BX1 i_1531927(
		.AN(n_1904),
		.B(op_a[24]),
		.C(op_a[25]),
		.D(n_2305),
		.Y(n_2372));

	OAI211X1 i_1435(
		.A0(op_a[26]),
		.A1(n_7313),
		.B0(op_b[26]),
		.C0(cmd[1]),
		.Y(n_2373));

	OAI221XL i_1437(
		.A0(n_1700),
		.A1(n_6901),
		.B0(n_1599),
		.B1(n_6911),
		.C0(n_2373),
		.Y(n_2375));

	AOI221X1 i_1439(
		.A0(n_6906),
		.A1(op_a[26]),
		.B0(n_1600),
		.B1(n_6904),
		.C0(n_2375),
		.Y(n_2377));

	OAI31X1 i_1440(
		.A0(n_2360),
		.A1(n_7323),
		.A2(n_1708),
		.B0(n_2377),
		.Y(n_2378));

	AOI21X1 i_271(
		.A0(op_a[27]),
		.A1(op_b[27]),
		.B0(n_1650),
		.Y(n_2382));

	OAI211X1 i_1465(
		.A0(op_a[27]),
		.A1(n_7313),
		.B0(op_b[27]),
		.C0(n_7320),
		.Y(n_2383));

	OAI21XL i_1466(
		.A0(n_1650),
		.A1(n_1942),
		.B0(n_2383),
		.Y(n_2384));

	AOI21X1 i_1467(
		.A0(n_7338),
		.A1(op_a[27]),
		.B0(n_2384),
		.Y(n_2385));

	OAI221XL i_1469(
		.A0(n_3068),
		.A1(n_1622),
		.B0(n_1623),
		.B1(n_3095),
		.C0(n_2385),
		.Y(n_2387));

	NOR2BX1 i_276(
		.AN(n_1706),
		.B(n_1710),
		.Y(n_2390));

	OAI2BB1X1 i_1887234(
		.A0N(n_1640),
		.A1N(n_1744),
		.B0(n_3069),
		.Y(n_2391));

	AOI31X1 i_440(
		.A0(n_1640),
		.A1(n_1709),
		.A2(n_1639),
		.B0(n_2391),
		.Y(n_2393));

	OAI211X1 i_1501(
		.A0(op_a[28]),
		.A1(n_7313),
		.B0(op_b[28]),
		.C0(n_7320),
		.Y(n_2394));

	OAI2BB1X1 i_1502(
		.A0N(n_3066),
		.A1N(n_3064),
		.B0(n_2394),
		.Y(n_2395));

	AOI211X1 i_1504(
		.A0(n_7338),
		.A1(op_a[28]),
		.B0(n_2395),
		.C0(n_1661),
		.Y(n_2397));

	OAI21XL i_1551509(
		.A0(n_1650),
		.A1(n_1817),
		.B0(n_1814),
		.Y(n_2399));

	NOR2BX1 i_403(
		.AN(n_1648),
		.B(n_2399),
		.Y(n_2401));

	AOI21X1 i_277(
		.A0(op_a[28]),
		.A1(op_b[28]),
		.B0(n_1697),
		.Y(n_2402));

	AOI32X1 i_1506(
		.A0(n_2393),
		.A1(n_3062),
		.A2(n_2390),
		.B0(n_1656),
		.B1(n_7341),
		.Y(n_2404));

	NAND2BX1 i_281(
		.AN(n_1713),
		.B(n_885),
		.Y(n_2406));

	OAI21XL i_1514(
		.A0(n_1750),
		.A1(n_3090),
		.B0(n_1746),
		.Y(n_2408));

	OAI21XL i_441(
		.A0(n_1670),
		.A1(n_1743),
		.B0(n_1742),
		.Y(n_2409));

	AOI21X1 i_1524(
		.A0(n_1823),
		.A1(n_3091),
		.B0(n_1819),
		.Y(n_2411));

	OAI21XL i_283(
		.A0(op_b[29]),
		.A1(op_a[29]),
		.B0(n_1812),
		.Y(n_2413));

	NOR4BX1 i_1561930(
		.AN(n_1908),
		.B(op_a[25]),
		.C(op_a[28]),
		.D(n_2352),
		.Y(n_2417));

	OAI211X1 i_1537(
		.A0(op_a[29]),
		.A1(n_7313),
		.B0(op_b[29]),
		.C0(n_7320),
		.Y(n_2418));

	OAI221XL i_1539(
		.A0(n_1703),
		.A1(n_1942),
		.B0(n_1682),
		.B1(n_3068),
		.C0(n_2418),
		.Y(n_2420));

	AOI211X1 i_1541(
		.A0(n_7338),
		.A1(op_a[29]),
		.B0(n_2420),
		.C0(n_1689),
		.Y(n_2422));

	OAI2BB1X1 i_1542(
		.A0N(n_1683),
		.A1N(n_7341),
		.B0(n_2422),
		.Y(n_2423));

	NAND2BX1 i_1587204(
		.AN(n_952),
		.B(n_954),
		.Y(n_2425));

	NOR2BX1 i_1565(
		.AN(n_1709),
		.B(n_1743),
		.Y(n_2426));

	OAI21XL i_442(
		.A0(n_1714),
		.A1(n_1713),
		.B0(n_885),
		.Y(n_2428));

	OAI21XL i_405(
		.A0(n_1704),
		.A1(n_1703),
		.B0(n_1812),
		.Y(n_2431));

	NAND3X1 i_1571931(
		.A(n_1912),
		.B(n_1908),
		.C(n_2372),
		.Y(n_2434));

	AOI211X1 i_1553(
		.A0(cmd[1]),
		.A1(op_b[30]),
		.B0(n_6906),
		.C0(n_3064),
		.Y(n_2436));

	NOR2BX1 i_1578(
		.AN(n_2434),
		.B(op_a[30]),
		.Y(n_2437));

	AOI222X1 i_1580(
		.A0(n_2437),
		.A1(n_1918),
		.B0(op_b[30]),
		.B1(n_1946),
		.C0(n_1720),
		.C1(op_a[30]),
		.Y(n_2439));

	OAI221XL i_1582(
		.A0(n_1915),
		.A1(n_3068),
		.B0(n_1723),
		.B1(n_2425),
		.C0(n_2439),
		.Y(n_2441));

	NOR4X1 i_81615(
		.A(cmd[0]),
		.B(cmd[2]),
		.C(cmd[3]),
		.D(cmd[1]),
		.Y(n_868));

	AOI21X1 i_1398(
		.A0(n_1738),
		.A1(n_3095),
		.B0(n_828),
		.Y(result[32]));

	NOR4BBX1 i_671598(
		.AN(n_1912),
		.BN(op_a[31]),
		.C(op_a[30]),
		.D(n_1911),
		.Y(n_166));

	NAND2X1 i_2154(
		.A(ovm),
		.B(result[32]),
		.Y(n_9076575));

	INVX1 i_3032(
		.A(n_827),
		.Y(n_3060));

	INVX1 i_3034(
		.A(n_1738),
		.Y(n_3062));

	INVX1 i_3035(
		.A(n_1944),
		.Y(n_3063));

	INVX1 i_3036(
		.A(n_6901),
		.Y(n_3064));

	INVX1 i_3037(
		.A(n_1136),
		.Y(n_3065));

	INVX1 i_3038(
		.A(n_1697),
		.Y(n_3066));

	INVX1 i_3039(
		.A(n_1886),
		.Y(n_3067));

	INVX1 i_3040(
		.A(n_1918),
		.Y(n_3068));

	INVX1 i_3041(
		.A(n_1741),
		.Y(n_3069));

	INVX1 i_3042(
		.A(n_1742),
		.Y(n_3070));

	INVX1 i_3043(
		.A(n_1808),
		.Y(n_3071));

	INVX1 i_3044(
		.A(n_984),
		.Y(result[0]));

	INVX1 i_3045(
		.A(n_1781),
		.Y(n_3073));

	INVX1 i_3046(
		.A(n_1784),
		.Y(n_3074));

	INVX1 i_3047(
		.A(n_1793),
		.Y(n_3075));

	INVX1 i_3048(
		.A(n_1213),
		.Y(n_3076));

	INVX1 i_3049(
		.A(n_1816),
		.Y(n_3077));

	INVX1 i_3050(
		.A(n_1853),
		.Y(n_3078));

	INVX1 i_3051(
		.A(n_1858),
		.Y(n_3079));

	INVX1 i_3052(
		.A(n_1857),
		.Y(n_3080));

	INVX1 i_3053(
		.A(n_1861),
		.Y(n_3081));

	INVX1 i_3054(
		.A(n_1860),
		.Y(n_3082));

	INVX1 i_3055(
		.A(n_1866),
		.Y(n_3083));

	INVX1 i_3056(
		.A(n_1865),
		.Y(n_3084));

	INVX1 i_3057(
		.A(n_1868),
		.Y(n_3085));

	INVX1 i_3058(
		.A(n_911),
		.Y(n_3086));

	INVX1 i_3059(
		.A(n_1996),
		.Y(n_3087));

	INVX1 i_3060(
		.A(n_2428),
		.Y(n_3088));

	INVX1 i_3061(
		.A(n_2040),
		.Y(n_3089));

	INVX1 i_3062(
		.A(n_2342),
		.Y(n_3090));

	INVX1 i_3063(
		.A(n_2346),
		.Y(n_3091));

	INVX1 i_3064(
		.A(n_2083),
		.Y(n_3092));

	INVX1 i_3065(
		.A(n_2344),
		.Y(n_3093));

	INVX1 i_3066(
		.A(n_9076575),
		.Y(n_907));

	INVX1 i_3067(
		.A(n_6904),
		.Y(n_3095));

endmodule
module data_bus_mach(
		clk,
		reset,
		read,
		write,
		address,
		data_in,
		data_out,
		pad_data_in,
		pad_data_out,
		addrs_in,
		read_cycle,
		sync,
		go,
		as,
		done,
		bus_request,
		bus_grant,
		scan_en,
		BG_scan_in,
		BG_scan_out,
	FE_PT1_,
	n_7867,
	FE_PT2_,
	SPCASCAN_N23_done,
	SPCASCAN_N24_t_sel_7,
	FE_PT3_,
	samp_bio,
	FE_PT4_);
   input FE_PT1_;
   input n_7867;
   input FE_PT2_;
   output SPCASCAN_N23_done;
   input SPCASCAN_N24_t_sel_7;
   input FE_PT3_;
   input samp_bio;
   input FE_PT4_;

	input clk;
	input reset;
	output read;
	output write;
	output [7:0] address;
	input [15:0] data_in;
	output [15:0] data_out;
	input [15:0] pad_data_in;
	output [15:0] pad_data_out;
	input [7:0] addrs_in;
	input read_cycle;
	input sync;
	input go;
	output as;
	output done;
	output bus_request;
	input bus_grant;
	input scan_en;
	input BG_scan_in;
	output BG_scan_out;

	wire [2:0] present_state;



	INVXL i_10642(
		.A(n_7893),
		.Y(BG_scan_out));

	INVXL i_10641(
		.A(bus_request),
		.Y(n_7893));

	CLKBUFXL i_10100(
		.A(n_4642),
		.Y(n_7173));

	CLKBUFX3 i_10050(
		.A(n_5177),
		.Y(n_7106));

	INVXL i_9590(
		.A(n_6389),
		.Y(pad_data_out[0]));

	INVXL i_9589(
		.A(data_in[0]),
		.Y(n_6389));

	BUFX3 i_9588(
		.A(data_in[1]),
		.Y(pad_data_out[1]));

	INVXL i_9584(
		.A(n_6381),
		.Y(pad_data_out[2]));

	INVXL i_9583(
		.A(data_in[2]),
		.Y(n_6381));

	CLKBUFX3 i_9582(
		.A(data_in[3]),
		.Y(pad_data_out[3]));

	INVXL i_9578(
		.A(n_6373),
		.Y(pad_data_out[4]));

	INVXL i_9577(
		.A(data_in[4]),
		.Y(n_6373));

	BUFX3 i_9576(
		.A(data_in[5]),
		.Y(pad_data_out[5]));

	BUFX3 i_9573(
		.A(data_in[6]),
		.Y(pad_data_out[6]));

	INVX1 i_9569(
		.A(n_6361),
		.Y(pad_data_out[8]));

	INVXL i_9568(
		.A(data_in[8]),
		.Y(n_6361));

	BUFX3 i_9567(
		.A(data_in[9]),
		.Y(pad_data_out[9]));

	INVXL i_9563(
		.A(n_6353),
		.Y(pad_data_out[10]));

	INVXL i_9562(
		.A(data_in[10]),
		.Y(n_6353));

	INVXL i_9560(
		.A(n_6349),
		.Y(pad_data_out[11]));

	INVXL i_9559(
		.A(data_in[11]),
		.Y(n_6349));

	CLKBUFX3 i_9558(
		.A(data_in[12]),
		.Y(pad_data_out[12]));

	INVXL i_9554(
		.A(n_6341),
		.Y(pad_data_out[13]));

	INVXL i_9553(
		.A(data_in[13]),
		.Y(n_6341));

	INVX1 i_9551(
		.A(n_6337),
		.Y(pad_data_out[14]));

	INVXL i_9550(
		.A(data_in[14]),
		.Y(n_6337));

	INVX1 i_9548(
		.A(n_6333),
		.Y(pad_data_out[15]));

	INVXL i_9547(
		.A(data_in[15]),
		.Y(n_6333));

	INVXL i_9545(
		.A(n_6329),
		.Y(address[1]));

	INVXL i_9544(
		.A(addrs_in[1]),
		.Y(n_6329));

	INVXL i_9542(
		.A(n_6325),
		.Y(address[4]));

	INVXL i_9541(
		.A(addrs_in[4]),
		.Y(n_6325));

	INVXL i_9539(
		.A(n_6321),
		.Y(address[5]));

	INVXL i_9538(
		.A(addrs_in[5]),
		.Y(n_6321));

	INVXL i_9536(
		.A(n_6317),
		.Y(address[6]));

	INVXL i_9535(
		.A(addrs_in[6]),
		.Y(n_6317));

	INVXL i_9533(
		.A(n_6313),
		.Y(address[7]));

	INVXL i_9532(
		.A(addrs_in[7]),
		.Y(n_6313));

	CLKBUFXL i_9491(
		.A(addrs_in[0]),
		.Y(address[0]));

	CLKBUFX3 i_9486(
		.A(addrs_in[3]),
		.Y(address[3]));

	CLKBUFX3 i_9485(
		.A(addrs_in[2]),
		.Y(address[2]));

	CLKBUFX3 i_9474(
		.A(data_in[7]),
		.Y(pad_data_out[7]));

	NOR2X1 i_11(
		.A(go),
		.B(present_state[2]),
		.Y(n_16));

	OAI21XL i_8(
		.A0(n_16),
		.A1(present_state[1]),
		.B0(n_23),
		.Y(n_21));

	SDFFRHQX1 present_state_reg_0(
		.SI(BG_scan_in),
		.SE(scan_en),
		.D(\nbus_626[0] ),
		.CK(clk),
		.RN(n_7173),
		.Q(present_state[0]));

	SDFFRHQX1 present_state_reg_1(
		.SI(data_out[15]),
		.SE(scan_en),
		.D(n_4641),
		.CK(clk),
		.RN(n_7173),
		.Q(present_state[1]));

	SDFFRHQX1 present_state_reg_2(
		.SI(FE_PT4_),
		.SE(scan_en),
		.D(n_24),
		.CK(clk),
		.RN(n_7173),
		.Q(present_state[2]));

	SDFFRHQX1 data_out_reg_0(
		.SI(data_out[7]),
		.SE(scan_en),
		.D(n_4534),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[0]));

	MX2X1 i_6145(
		.S0(n_7106),
		.B(pad_data_in[0]),
		.A(data_out[0]),
		.Y(n_4534));

	SDFFRHQX1 data_out_reg_1(
		.SI(FE_PT2_),
		.SE(scan_en),
		.D(n_4540),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[1]));

	MX2X1 i_6152(
		.S0(n_7106),
		.B(pad_data_in[1]),
		.A(data_out[1]),
		.Y(n_4540));

	XNOR2X1 i_3(
		.A(present_state[0]),
		.B(present_state[1]),
		.Y(n_23));

	SDFFRHQX1 data_out_reg_2(
		.SI(FE_PT1_),
		.SE(scan_en),
		.D(n_4546),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[2]));

	MX2X1 i_6159(
		.S0(n_7106),
		.B(pad_data_in[2]),
		.A(data_out[2]),
		.Y(n_4546));

	OAI32X1 i_2(
		.A0(present_state[1]),
		.A1(present_state[0]),
		.A2(n_28),
		.B0(n_5205),
		.B1(n_4640),
		.Y(n_24));

	SDFFRHQX1 data_out_reg_3(
		.SI(data_out[2]),
		.SE(scan_en),
		.D(n_4552),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[3]));

	MX2X1 i_6166(
		.S0(n_7106),
		.B(pad_data_in[3]),
		.A(data_out[3]),
		.Y(n_4552));

	SDFFRHQX1 data_out_reg_4(
		.SI(data_out[6]),
		.SE(scan_en),
		.D(n_4558),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[4]));

	MX2X1 i_6173(
		.S0(n_7106),
		.B(pad_data_in[4]),
		.A(data_out[4]),
		.Y(n_4558));

	SDFFRHQX1 data_out_reg_5(
		.SI(n_7867),
		.SE(scan_en),
		.D(n_4564),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[5]));

	MX2X1 i_6180(
		.S0(n_7106),
		.B(pad_data_in[5]),
		.A(data_out[5]),
		.Y(n_4564));

	SDFFRHQX1 data_out_reg_6(
		.SI(data_out[3]),
		.SE(scan_en),
		.D(n_4570),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[6]));

	MX2X1 i_6187(
		.S0(n_7106),
		.B(pad_data_in[6]),
		.A(data_out[6]),
		.Y(n_4570));

	NAND3BX1 i_26(
		.AN(read_cycle),
		.B(bus_grant),
		.C(go),
		.Y(n_28));

	SDFFRHQX1 data_out_reg_7(
		.SI(data_out[5]),
		.SE(scan_en),
		.D(n_4576),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[7]));

	MX2X1 i_6194(
		.S0(n_7106),
		.B(pad_data_in[7]),
		.A(data_out[7]),
		.Y(n_4576));

	SDFFRHQX1 data_out_reg_8(
		.SI(SPCASCAN_N24_t_sel_7),
		.SE(scan_en),
		.D(n_4582),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[8]));

	MX2X1 i_6201(
		.S0(n_7106),
		.B(pad_data_in[8]),
		.A(data_out[8]),
		.Y(n_4582));

	SDFFRHQX1 data_out_reg_9(
		.SI(data_out[13]),
		.SE(scan_en),
		.D(n_4588),
		.CK(clk),
		.RN(n_4642),
		.Q(data_out[9]));

	MX2X1 i_6208(
		.S0(n_7106),
		.B(pad_data_in[9]),
		.A(data_out[9]),
		.Y(n_4588));

	AOI31X1 i_20(
		.A0(bus_grant),
		.A1(read_cycle),
		.A2(go),
		.B0(present_state[1]),
		.Y(n_31));

	SDFFRHQX1 data_out_reg_10(
		.SI(as),
		.SE(scan_en),
		.D(n_4594),
		.CK(clk),
		.RN(n_4642),
		.Q(data_out[10]));

	MX2X1 i_6215(
		.S0(n_5177),
		.B(pad_data_in[10]),
		.A(data_out[10]),
		.Y(n_4594));

	SDFFRHQX1 data_out_reg_11(
		.SI(present_state[0]),
		.SE(scan_en),
		.D(n_4600),
		.CK(clk),
		.RN(n_4642),
		.Q(data_out[11]));

	MX2X1 i_6222(
		.S0(n_7106),
		.B(pad_data_in[11]),
		.A(data_out[11]),
		.Y(n_4600));

	NOR3X1 i_0(
		.A(present_state[0]),
		.B(present_state[1]),
		.C(n_4640),
		.Y(n_5232));

	SDFFRHQX1 data_out_reg_12(
		.SI(data_out[9]),
		.SE(scan_en),
		.D(n_4606),
		.CK(clk),
		.RN(n_4642),
		.Q(data_out[12]));

	MX2X1 i_6229(
		.S0(n_7106),
		.B(pad_data_in[12]),
		.A(data_out[12]),
		.Y(n_4606));

	NOR3BX1 i_19008(
		.AN(present_state[0]),
		.B(present_state[1]),
		.C(present_state[2]),
		.Y(n_5226));

	SDFFRHQX1 data_out_reg_13(
		.SI(data_out[14]),
		.SE(scan_en),
		.D(n_4612),
		.CK(clk),
		.RN(n_4642),
		.Q(data_out[13]));

	MX2X1 i_6236(
		.S0(n_7106),
		.B(pad_data_in[13]),
		.A(data_out[13]),
		.Y(n_4612));

	AOI21X1 i_5(
		.A0(n_31),
		.A1(n_4640),
		.B0(present_state[0]),
		.Y(\nbus_626[0] ));

	SDFFRHQX1 data_out_reg_14(
		.SI(FE_PT3_),
		.SE(scan_en),
		.D(n_4618),
		.CK(clk),
		.RN(n_4642),
		.Q(data_out[14]));

	MX2X1 i_6243(
		.S0(n_7106),
		.B(pad_data_in[14]),
		.A(data_out[14]),
		.Y(n_4618));

	AND2X1 i_7(
		.A(present_state[0]),
		.B(present_state[1]),
		.Y(n_5205));

	SDFFRHQX1 data_out_reg_15(
		.SI(data_out[8]),
		.SE(scan_en),
		.D(n_4624),
		.CK(clk),
		.RN(n_7173),
		.Q(data_out[15]));

	MX2X1 i_6250(
		.S0(n_7106),
		.B(pad_data_in[15]),
		.A(data_out[15]),
		.Y(n_4624));

	NOR3BX1 i_9(
		.AN(present_state[1]),
		.B(present_state[0]),
		.C(present_state[2]),
		.Y(n_5177));

	DFFRHQX1 write_reg(
		.D(n_5232),
		.CK(clk),
		.RN(n_4642),
		.Q(write));

	SDFFRHQX1 read_reg(
		.SI(present_state[2]),
		.SE(scan_en),
		.D(n_5226),
		.CK(clk),
		.RN(n_7173),
		.Q(read));

	SDFFRHQX1 done_reg(
		.SI(present_state[1]),
		.SE(scan_en),
		.D(n_5205),
		.CK(clk),
		.RN(n_7173),
		.Q(SPCASCAN_N23_done));

	SDFFRHQX1 as_reg(
		.SI(BG_scan_out),
		.SE(scan_en),
		.D(n_21),
		.CK(clk),
		.RN(n_4642),
		.Q(as));

	SDFFRHQX1 bus_request_reg(
		.SI(samp_bio),
		.SE(scan_en),
		.D(n_21),
		.CK(clk),
		.RN(n_4642),
		.Q(bus_request));

	INVX1 i_6322(
		.A(present_state[2]),
		.Y(n_4640));

	INVX1 i_6323(
		.A(n_23),
		.Y(n_4641));

	INVX1 i_6324(
		.A(reset),
		.Y(n_4642));

endmodule
module decode_i(
		clk,
		reset,
		phi_1,
		phi_2,
		phi_3,
		phi_4,
		phi_5,
		phi_6,
		decode,
		p_data_out,
		ir,
		skip_one,
		read_prog,
		go_prog,
		read_data,
		go_data,
		read_port,
		go_port,
		decode_skip_one,
		scan_en,
		BG_scan_in,
		BG_scan_out,
	FE_PT1_,
	FE_PT2_,
	FE_PT3_,
	FE_PT4_,
	FE_PT5_,
	FE_PT6_,
	FE_PT7_,
	FE_PT8_,
	arp,
	pc_acc,
	SPCASCAN_N34_two_cycle,
	enc_read_port,
	UNCONNECTED_006,
	enc_go_data,
	enc_read_data);
   input FE_PT1_;
   input FE_PT2_;
   input FE_PT3_;
   input FE_PT4_;
   input FE_PT5_;
   input FE_PT6_;
   input FE_PT7_;
   input FE_PT8_;
   input arp;
   input pc_acc;
   output SPCASCAN_N34_two_cycle;
   input enc_read_port;
   input UNCONNECTED_006;
   input enc_go_data;
   input enc_read_data;

	input clk;
	input reset;
	input phi_1;
	input phi_2;
	input phi_3;
	input phi_4;
	input phi_5;
	input phi_6;
	output [15:0] decode;
	input [15:0] p_data_out;
	output [15:0] ir;
	input skip_one;
	output read_prog;
	output go_prog;
	output read_data;
	output go_data;
	output read_port;
	output go_port;
	output decode_skip_one;
	input scan_en;
	input BG_scan_in;
	output BG_scan_out;




	CLKBUFXL i_10129(
		.A(n_4475),
		.Y(n_7215));

	CLKBUFXL i_10126(
		.A(n_7043),
		.Y(n_7212));

	CLKBUFX3 i_10108(
		.A(n_4475),
		.Y(n_7185));

	BUFX1 i_10107(
		.A(n_181),
		.Y(n_7182));

	CLKBUFXL i_10028(
		.A(\nbus_708[15] ),
		.Y(ir[15]));

	CLKBUFX3 i_10013(
		.A(n_181),
		.Y(n_7043));

	CLKBUFXL i_9919(
		.A(\nbus_669[15] ),
		.Y(decode[15]));

	BUFX3 i_9918(
		.A(decode[11]),
		.Y(n_7361));

	BUFX3 i_9917(
		.A(decode[12]),
		.Y(n_7366));

	OAI21XL i_58(
		.A0(n_73),
		.A1(n_140),
		.B0(n_4472),
		.Y(n_74));

	NOR3X1 i_56(
		.A(decode[12]),
		.B(n_129),
		.C(n_143),
		.Y(n_73));

	NOR2BX1 i_1036(
		.AN(n_179),
		.B(phi_3),
		.Y(n_438));

	NOR2BX1 i_947(
		.AN(n_753),
		.B(phi_3),
		.Y(n_408));

	AND2X1 i_574(
		.A(n_68),
		.B(n_124),
		.Y(n_753));

	NAND4X1 i_35(
		.A(n_123),
		.B(n_122),
		.C(n_107),
		.D(n_176),
		.Y(n_69));

	NAND2BX1 i_33(
		.AN(n_181),
		.B(decode_skip_one),
		.Y(n_68));

	NAND2X1 i_61(
		.A(decode[9]),
		.B(n_152),
		.Y(n_75));

	NAND3X1 i_62(
		.A(decode[8]),
		.B(decode[10]),
		.C(decode[11]),
		.Y(n_76));

	NAND3X1 i_36(
		.A(n_132),
		.B(n_76),
		.C(n_75),
		.Y(n_79));

	OAI21XL i_27(
		.A0(decode[9]),
		.A1(n_146),
		.B0(n_7366),
		.Y(n_82));

	OAI21XL i_40(
		.A0(decode[8]),
		.A1(decode[11]),
		.B0(n_118),
		.Y(n_83));

	AOI211X1 i_74(
		.A0(decode[13]),
		.A1(n_4473),
		.B0(decode[14]),
		.C0(decode[15]),
		.Y(n_84));

	NAND3X1 i_79(
		.A(n_150),
		.B(n_161),
		.C(n_135),
		.Y(n_88));

	NOR4X1 i_82(
		.A(decode[10]),
		.B(decode[11]),
		.C(decode[9]),
		.D(n_145),
		.Y(n_90));

	NAND4BBX1 i_34(
		.AN(n_139),
		.BN(n_163),
		.C(n_165),
		.D(n_134),
		.Y(n_92));

	AOI21X1 i_1009(
		.A0(n_92),
		.A1(n_4472),
		.B0(phi_3),
		.Y(n_564));

	AOI22X1 i_25(
		.A0(decode[10]),
		.A1(n_141),
		.B0(decode[11]),
		.B1(n_4471),
		.Y(n_95));

	OAI21XL i_808(
		.A0(n_95),
		.A1(n_169),
		.B0(n_68),
		.Y(n_576));

	OAI21XL i_570(
		.A0(n_165),
		.A1(n_124),
		.B0(n_183),
		.Y(n_831));

	NAND2X1 i_24(
		.A(decode[11]),
		.B(n_130),
		.Y(n_99));

	OAI2BB1X1 i_31(
		.A0N(decode[14]),
		.A1N(n_99),
		.B0(decode[13]),
		.Y(n_101));

	NOR2X1 i_99(
		.A(n_139),
		.B(decode[15]),
		.Y(n_102));

	AOI221X1 i_38(
		.A0(decode[14]),
		.A1(n_132),
		.B0(decode[15]),
		.B1(n_101),
		.C0(n_102),
		.Y(n_105));

	OAI21XL i_630(
		.A0(n_105),
		.A1(n_124),
		.B0(n_68),
		.Y(n_411));

	NAND3BX1 i_107(
		.AN(n_133),
		.B(n_130),
		.C(n_143),
		.Y(n_107));

	NOR2X1 i_111(
		.A(decode[10]),
		.B(n_4471),
		.Y(n_109));

	AOI21X1 i_112(
		.A0(decode[10]),
		.A1(n_141),
		.B0(decode[11]),
		.Y(n_110));

	NOR2BX1 i_113(
		.AN(n_148),
		.B(n_156),
		.Y(n_112));

	AOI2BB1X1 i_114(
		.A0N(n_110),
		.A1N(n_109),
		.B0(n_129),
		.Y(n_113));

	AOI21X1 i_28(
		.A0(n_146),
		.A1(n_149),
		.B0(decode[9]),
		.Y(n_115));

	AOI31X1 i_30(
		.A0(n_150),
		.A1(n_161),
		.A2(decode[14]),
		.B0(decode[13]),
		.Y(n_116));

	NAND2BX1 i_18(
		.AN(n_149),
		.B(decode[9]),
		.Y(n_118));

	NAND2X1 i_118(
		.A(decode[15]),
		.B(n_116),
		.Y(n_122));

	OAI21XL i_119(
		.A0(n_113),
		.A1(n_112),
		.B0(decode[12]),
		.Y(n_123));

	NAND2BX1 i_09006(
		.AN(n_181),
		.B(n_182),
		.Y(n_124));

	NOR2BX1 i_23(
		.AN(decode[13]),
		.B(decode[14]),
		.Y(n_125));

	NAND2X1 i_46(
		.A(decode[14]),
		.B(decode[13]),
		.Y(n_128));

	NAND3X1 i_277(
		.A(decode[14]),
		.B(decode[13]),
		.C(decode[15]),
		.Y(n_129));

	NOR2X1 i_346(
		.A(decode[12]),
		.B(n_129),
		.Y(n_130));

	NAND3BX1 i_3(
		.AN(decode[9]),
		.B(decode[8]),
		.C(decode[10]),
		.Y(n_132));

	NOR2BX1 i_17(
		.AN(decode[11]),
		.B(n_132),
		.Y(n_133));

	AOI32X1 i_1(
		.A0(decode[15]),
		.A1(n_125),
		.A2(decode[12]),
		.B0(n_130),
		.B1(n_133),
		.Y(n_134));

	NOR2BX1 i_4(
		.AN(decode[14]),
		.B(decode[13]),
		.Y(n_135));

	NOR4BX1 i_281(
		.AN(decode[14]),
		.B(decode[15]),
		.C(n_7366),
		.D(decode[13]),
		.Y(n_137));

	NOR3BX1 i_292(
		.AN(n_137),
		.B(n_132),
		.C(decode[11]),
		.Y(n_139));

	NAND2BX1 i_12(
		.AN(n_139),
		.B(n_134),
		.Y(n_140));

	NAND2X1 i_8(
		.A(decode[8]),
		.B(decode[9]),
		.Y(n_141));

	SDFFRHQX1 two_cycle_reg(
		.SI(read_port),
		.SE(scan_en),
		.D(n_4225),
		.CK(clk),
		.RN(n_7215),
		.Q(SPCASCAN_N34_two_cycle));

	OAI211X1 i_5212(
		.A0(n_179),
		.A1(n_438),
		.B0(n_74),
		.C0(n_4228),
		.Y(n_4225));

	NAND3X1 i_5214(
		.A(n_74),
		.B(n_438),
		.C(SPCASCAN_N34_two_cycle),
		.Y(n_4228));

	NAND4BXL i_48(
		.AN(decode[11]),
		.B(decode[10]),
		.C(decode[8]),
		.D(decode[9]),
		.Y(n_143));

	SDFFRHQX1 decode_skip_one_reg(
		.SI(enc_read_data),
		.SE(scan_en),
		.D(n_4231),
		.CK(clk),
		.RN(n_7215),
		.Q(decode_skip_one));

	MX2X1 i_5219(
		.S0(n_576),
		.B(n_182),
		.A(decode_skip_one),
		.Y(n_4231));

	NOR2BX1 i_67(
		.AN(decode[12]),
		.B(decode[15]),
		.Y(n_144));

	SDFFRHQX1 decode_reg_0(
		.SI(decode[5]),
		.SE(scan_en),
		.D(n_4237),
		.CK(clk),
		.RN(n_7215),
		.Q(decode[0]));

	MX2X1 i_5226(
		.S0(n_7043),
		.B(decode[0]),
		.A(p_data_out[0]),
		.Y(n_4237));

	NAND2X1 i_422(
		.A(n_125),
		.B(n_144),
		.Y(n_145));

	SDFFRHQX1 decode_reg_1(
		.SI(FE_PT7_),
		.SE(scan_en),
		.D(n_4243),
		.CK(clk),
		.RN(n_7215),
		.Q(decode[1]));

	MX2X1 i_5233(
		.S0(n_7043),
		.B(decode[1]),
		.A(p_data_out[1]),
		.Y(n_4243));

	NAND2BX1 i_11(
		.AN(decode[10]),
		.B(n_7361),
		.Y(n_146));

	SDFFRHQX1 decode_reg_2(
		.SI(decode[0]),
		.SE(scan_en),
		.D(n_4249),
		.CK(clk),
		.RN(n_7215),
		.Q(decode[2]));

	MX2X1 i_5240(
		.S0(n_7043),
		.B(decode[2]),
		.A(p_data_out[2]),
		.Y(n_4249));

	SDFFRHQX1 decode_reg_3(
		.SI(ir[5]),
		.SE(scan_en),
		.D(n_4255),
		.CK(clk),
		.RN(n_4475),
		.Q(decode[3]));

	MX2X1 i_5247(
		.S0(n_7043),
		.B(decode[3]),
		.A(p_data_out[3]),
		.Y(n_4255));

	NOR2X1 i_269(
		.A(decode[15]),
		.B(n_128),
		.Y(n_148));

	SDFFRHQX1 decode_reg_4(
		.SI(FE_PT6_),
		.SE(scan_en),
		.D(n_4261),
		.CK(clk),
		.RN(n_7215),
		.Q(decode[4]));

	MX2X1 i_5254(
		.S0(n_7043),
		.B(decode[4]),
		.A(p_data_out[4]),
		.Y(n_4261));

	OR2X1 i_5(
		.A(decode[10]),
		.B(n_7361),
		.Y(n_149));

	SDFFRHQX1 decode_reg_5(
		.SI(FE_PT4_),
		.SE(scan_en),
		.D(n_4267),
		.CK(clk),
		.RN(n_7215),
		.Q(decode[5]));

	MX2X1 i_5261(
		.S0(n_7043),
		.B(decode[5]),
		.A(p_data_out[5]),
		.Y(n_4267));

	NOR2X1 i_15(
		.A(n_7366),
		.B(n_149),
		.Y(n_150));

	SDFFRHQX1 decode_reg_6(
		.SI(FE_PT5_),
		.SE(scan_en),
		.D(n_4273),
		.CK(clk),
		.RN(n_7215),
		.Q(decode[6]));

	MX2X1 i_5268(
		.S0(n_7043),
		.B(decode[6]),
		.A(p_data_out[6]),
		.Y(n_4273));

	NOR2BX1 i_22(
		.AN(n_148),
		.B(n_7366),
		.Y(n_151));

	SDFFSHQX1 decode_reg_7(
		.SI(ir[7]),
		.SE(scan_en),
		.D(n_4279),
		.CK(clk),
		.SN(n_7185),
		.Q(decode[7]));

	MX2X1 i_5275(
		.S0(n_7182),
		.B(decode[7]),
		.A(p_data_out[7]),
		.Y(n_4279));

	NOR2X1 i_10(
		.A(decode[8]),
		.B(n_7361),
		.Y(n_152));

	SDFFSHQX1 decode_reg_8(
		.SI(BG_scan_in),
		.SE(scan_en),
		.D(n_4285),
		.CK(clk),
		.SN(n_7185),
		.Q(decode[8]));

	MX2X1 i_5282(
		.S0(n_7182),
		.B(decode[8]),
		.A(p_data_out[8]),
		.Y(n_4285));

	SDFFSHQX1 decode_reg_9(
		.SI(decode[10]),
		.SE(scan_en),
		.D(n_4291),
		.CK(clk),
		.SN(n_7185),
		.Q(decode[9]));

	MX2X1 i_5289(
		.S0(n_7043),
		.B(decode[9]),
		.A(p_data_out[9]),
		.Y(n_4291));

	SDFFSHQX1 decode_reg_10(
		.SI(ir[11]),
		.SE(scan_en),
		.D(n_4297),
		.CK(clk),
		.SN(n_7185),
		.Q(decode[10]));

	MX2X1 i_5296(
		.S0(n_7182),
		.B(decode[10]),
		.A(p_data_out[10]),
		.Y(n_4297));

	AOI22X1 i_515(
		.A0(n_151),
		.A1(n_79),
		.B0(n_148),
		.B1(n_150),
		.Y(n_155));

	SDFFSHQX1 decode_reg_11(
		.SI(FE_PT2_),
		.SE(scan_en),
		.D(n_4303),
		.CK(clk),
		.SN(n_7185),
		.Q(decode[11]));

	MX2X1 i_5303(
		.S0(n_7182),
		.B(decode[11]),
		.A(p_data_out[11]),
		.Y(n_4303));

	AOI21X1 i_20(
		.A0(decode[8]),
		.A1(decode[9]),
		.B0(n_146),
		.Y(n_156));

	SDFFSHQX1 decode_reg_12(
		.SI(decode[1]),
		.SE(scan_en),
		.D(n_4309),
		.CK(clk),
		.SN(n_4475),
		.Q(decode[12]));

	MX2X1 i_5310(
		.S0(n_7182),
		.B(decode[12]),
		.A(p_data_out[12]),
		.Y(n_4309));

	SDFFSHQX1 decode_reg_13(
		.SI(FE_PT1_),
		.SE(scan_en),
		.D(n_4315),
		.CK(clk),
		.SN(n_7185),
		.Q(decode[13]));

	MX2X1 i_5317(
		.S0(n_7182),
		.B(decode[13]),
		.A(p_data_out[13]),
		.Y(n_4315));

	AOI32X1 i_77(
		.A0(decode[12]),
		.A1(n_148),
		.A2(n_156),
		.B0(n_137),
		.B1(n_83),
		.Y(n_158));

	SDFFSHQX1 decode_reg_14(
		.SI(ir[9]),
		.SE(scan_en),
		.D(n_4321),
		.CK(clk),
		.SN(n_7185),
		.Q(decode[14]));

	MX2X1 i_5324(
		.S0(n_7182),
		.B(decode[14]),
		.A(p_data_out[14]),
		.Y(n_4321));

	SDFFRHQX1 decode_reg_15(
		.SI(decode[11]),
		.SE(scan_en),
		.D(n_4327),
		.CK(clk),
		.RN(n_7215),
		.Q(\nbus_669[15] ));

	MX2X1 i_5331(
		.S0(n_7043),
		.B(decode[15]),
		.A(p_data_out[15]),
		.Y(n_4327));

	SDFFRHQX1 go_port_reg(
		.SI(pc_acc),
		.SE(scan_en),
		.D(n_4333),
		.CK(clk),
		.RN(n_7215),
		.Q(go_port));

	OAI21XL i_5338(
		.A0(n_179),
		.A1(n_438),
		.B0(n_4336),
		.Y(n_4333));

	NAND2X1 i_5340(
		.A(n_438),
		.B(go_port),
		.Y(n_4336));

	NOR2X1 i_9(
		.A(decode[8]),
		.B(decode[9]),
		.Y(n_161));

	SDFFRHQX1 go_data_reg(
		.SI(enc_go_data),
		.SE(scan_en),
		.D(n_4339),
		.CK(clk),
		.RN(n_7215),
		.Q(go_data));

	OAI2BB1X1 i_5345(
		.A0N(n_564),
		.A1N(go_data),
		.B0(n_4341),
		.Y(n_4339));

	NAND2BX1 i_5346(
		.AN(n_564),
		.B(n_831),
		.Y(n_4341));

	SDFFRHQX1 read_prog_reg(
		.SI(BG_scan_out),
		.SE(scan_en),
		.D(n_4345),
		.CK(clk),
		.RN(n_7215),
		.Q(read_prog));

	OAI21XL i_5352(
		.A0(n_753),
		.A1(n_408),
		.B0(n_4348),
		.Y(n_4345));

	NAND2X1 i_5354(
		.A(n_408),
		.B(read_prog),
		.Y(n_4348));

	NAND4BXL i_13(
		.AN(n_84),
		.B(n_158),
		.C(n_155),
		.D(n_88),
		.Y(n_163));

	SDFFRHQX1 ir_reg_0(
		.SI(FE_PT3_),
		.SE(scan_en),
		.D(n_4351),
		.CK(clk),
		.RN(n_7215),
		.Q(ir[0]));

	MX2X1 i_5359(
		.S0(n_7043),
		.B(ir[0]),
		.A(decode[0]),
		.Y(n_4351));

	SDFFRHQX1 ir_reg_1(
		.SI(FE_PT8_),
		.SE(scan_en),
		.D(n_4357),
		.CK(clk),
		.RN(n_7215),
		.Q(ir[1]));

	MX2X1 i_5366(
		.S0(n_7043),
		.B(ir[1]),
		.A(decode[1]),
		.Y(n_4357));

	AOI21X1 i_14(
		.A0(n_135),
		.A1(n_144),
		.B0(n_90),
		.Y(n_165));

	SDFFRHQX1 ir_reg_2(
		.SI(ir[3]),
		.SE(scan_en),
		.D(n_4363),
		.CK(clk),
		.RN(n_7215),
		.Q(ir[2]));

	MX2X1 i_5373(
		.S0(n_7043),
		.B(ir[2]),
		.A(decode[2]),
		.Y(n_4363));

	SDFFRHQX1 ir_reg_3(
		.SI(ir[0]),
		.SE(scan_en),
		.D(n_4369),
		.CK(clk),
		.RN(n_4475),
		.Q(ir[3]));

	MX2X1 i_5380(
		.S0(n_7212),
		.B(ir[3]),
		.A(decode[3]),
		.Y(n_4369));

	SDFFRHQX1 ir_reg_4(
		.SI(decode[3]),
		.SE(scan_en),
		.D(n_4375),
		.CK(clk),
		.RN(n_4475),
		.Q(ir[4]));

	MX2X1 i_5387(
		.S0(n_7212),
		.B(ir[4]),
		.A(decode[4]),
		.Y(n_4375));

	SDFFRHQX1 ir_reg_5(
		.SI(decode[7]),
		.SE(scan_en),
		.D(n_4381),
		.CK(clk),
		.RN(n_4475),
		.Q(ir[5]));

	MX2X1 i_5394(
		.S0(n_7043),
		.B(ir[5]),
		.A(decode[5]),
		.Y(n_4381));

	NAND3BX1 i_92(
		.AN(n_129),
		.B(decode[12]),
		.C(n_4472),
		.Y(n_169));

	SDFFRHQX1 ir_reg_6(
		.SI(ir[4]),
		.SE(scan_en),
		.D(n_4387),
		.CK(clk),
		.RN(n_4475),
		.Q(ir[6]));

	MX2X1 i_5401(
		.S0(n_7212),
		.B(ir[6]),
		.A(decode[6]),
		.Y(n_4387));

	SDFFSHQX1 ir_reg_7(
		.SI(decode[12]),
		.SE(scan_en),
		.D(n_4393),
		.CK(clk),
		.SN(n_7185),
		.Q(ir[7]));

	MX2X1 i_5408(
		.S0(n_7182),
		.B(ir[7]),
		.A(decode[7]),
		.Y(n_4393));

	SDFFSHQX1 ir_reg_8(
		.SI(\nbus_669[15] ),
		.SE(scan_en),
		.D(n_4399),
		.CK(clk),
		.SN(n_7185),
		.Q(ir[8]));

	MX2X1 i_5415(
		.S0(n_7182),
		.B(ir[8]),
		.A(decode[8]),
		.Y(n_4399));

	SDFFSHQX1 ir_reg_9(
		.SI(ir[14]),
		.SE(scan_en),
		.D(n_4405),
		.CK(clk),
		.SN(n_7185),
		.Q(ir[9]));

	MX2X1 i_5422(
		.S0(n_7182),
		.B(ir[9]),
		.A(decode[9]),
		.Y(n_4405));

	SDFFSHQX1 ir_reg_10(
		.SI(arp),
		.SE(scan_en),
		.D(n_4411),
		.CK(clk),
		.SN(n_7185),
		.Q(ir[10]));

	MX2X1 i_5429(
		.S0(n_7182),
		.B(ir[10]),
		.A(decode[10]),
		.Y(n_4411));

	OAI211X1 i_122(
		.A0(decode[8]),
		.A1(decode[11]),
		.B0(n_137),
		.C0(n_118),
		.Y(n_174));

	SDFFSHQX1 ir_reg_11(
		.SI(\nbus_708[15] ),
		.SE(scan_en),
		.D(n_4417),
		.CK(clk),
		.SN(n_7185),
		.Q(ir[11]));

	MX2X1 i_5436(
		.S0(n_7182),
		.B(ir[11]),
		.A(decode[11]),
		.Y(n_4417));

	OAI22X1 i_123(
		.A0(n_139),
		.A1(n_174),
		.B0(n_115),
		.B1(n_145),
		.Y(n_175));

	SDFFSHQX1 ir_reg_12(
		.SI(decode[9]),
		.SE(scan_en),
		.D(n_4423),
		.CK(clk),
		.SN(n_7185),
		.Q(ir[12]));

	MX2X1 i_5443(
		.S0(n_7182),
		.B(ir[12]),
		.A(decode[12]),
		.Y(n_4423));

	AOI21X1 i_124(
		.A0(n_151),
		.A1(n_155),
		.B0(n_175),
		.Y(n_176));

	SDFFSHQX1 ir_reg_13(
		.SI(ir[10]),
		.SE(scan_en),
		.D(n_4429),
		.CK(clk),
		.SN(n_7185),
		.Q(ir[13]));

	MX2X1 i_5450(
		.S0(n_7182),
		.B(ir[13]),
		.A(decode[13]),
		.Y(n_4429));

	SDFFSHQX1 ir_reg_14(
		.SI(ir[13]),
		.SE(scan_en),
		.D(n_4435),
		.CK(clk),
		.SN(n_7185),
		.Q(ir[14]));

	MX2X1 i_5457(
		.S0(n_7182),
		.B(ir[14]),
		.A(decode[14]),
		.Y(n_4435));

	SDFFRHQX1 ir_reg_15(
		.SI(decode[14]),
		.SE(scan_en),
		.D(n_4441),
		.CK(clk),
		.RN(n_4475),
		.Q(\nbus_708[15] ));

	MX2X1 i_5464(
		.S0(n_7043),
		.B(ir[15]),
		.A(decode[15]),
		.Y(n_4441));

	NAND4BXL i_401(
		.AN(decode[12]),
		.B(decode[15]),
		.C(n_125),
		.D(n_4472),
		.Y(n_179));

	SDFFRHQX1 read_data_reg(
		.SI(UNCONNECTED_006),
		.SE(scan_en),
		.D(n_4447),
		.CK(clk),
		.RN(n_4475),
		.Q(read_data));

	OAI21XL i_5471(
		.A0(n_183),
		.A1(n_564),
		.B0(n_4450),
		.Y(n_4447));

	NAND2X1 i_5473(
		.A(n_564),
		.B(read_data),
		.Y(n_4450));

	NAND3BX1 i_663(
		.AN(n_124),
		.B(n_69),
		.C(n_4475),
		.Y(n_180));

	SDFFRHQX1 read_port_reg(
		.SI(enc_read_port),
		.SE(scan_en),
		.D(n_4453),
		.CK(clk),
		.RN(n_4475),
		.Q(read_port));

	OAI21XL i_5478(
		.A0(n_179),
		.A1(n_438),
		.B0(n_4456),
		.Y(n_4453));

	NAND2X1 i_5480(
		.A(n_438),
		.B(read_port),
		.Y(n_4456));

	NAND2BX1 i_2(
		.AN(skip_one),
		.B(phi_6),
		.Y(n_181));

	SDFFRHQX1 go_prog_reg(
		.SI(read_prog),
		.SE(scan_en),
		.D(n_4474),
		.CK(clk),
		.RN(n_4475),
		.Q(go_prog));

	AOI21X1 i_5485(
		.A0(n_408),
		.A1(go_prog),
		.B0(n_4461),
		.Y(n_4459));

	NOR2BX1 i_5486(
		.AN(n_411),
		.B(n_408),
		.Y(n_4461));

	NOR2X1 i_21123(
		.A(decode_skip_one),
		.B(SPCASCAN_N34_two_cycle),
		.Y(n_182));

	SDFFHQX1 null_op_reg(
		.SI(decode_skip_one),
		.SE(scan_en),
		.D(n_4468),
		.CK(clk),
		.Q(BG_scan_out));

	AND2X1 i_5494(
		.A(n_180),
		.B(BG_scan_out),
		.Y(n_4468));

	OAI21XL i_615(
		.A0(n_140),
		.A1(n_163),
		.B0(n_4472),
		.Y(n_183));

	INVX1 i_5659(
		.A(n_161),
		.Y(n_4471));

	INVX1 i_5660(
		.A(n_124),
		.Y(n_4472));

	INVX1 i_5661(
		.A(n_82),
		.Y(n_4473));

	INVX1 i_5662(
		.A(n_4459),
		.Y(n_4474));

	INVX1 i_5663(
		.A(reset),
		.Y(n_4475));

endmodule
module execute_i(
		clk,
		reset,
		phi_1,
		phi_2,
		phi_3,
		phi_4,
		phi_5,
		phi_6,
		decode_skip_one,
		gez,
		gz,
		nz,
		z,
		lz,
		lez,
		ov,
		arnz,
		bioz,
		alu_result,
		mpy_result,
		mdr,
		pdr,
		ir,
		decode,
		ar,
		skip_one,
		fetch_branch,
		branch_stall,
		pc_acc,
		dmov_inc,
		dp,
		arp,
		ar0,
		ar1,
		pc,
		acc,
		p,
		top,
		alu_cmd,
		sel_op_a,
		sel_op_b,
		read_prog,
		go_prog,
		read_data,
		go_data,
		read_port,
		go_port,
		ovm,
		scan_en,
		BG_scan_in,
		BG_scan_out,
	SPCASCAN_N6_present_state_2_,
	SPCASCAN_N7_present_state_1_,
	FE_PT1_,
	SPCASCAN_N23_done,
	SPCASCAN_N28_read,
	port_as,
	FE_PT2_,
	dec_go_port,
	SPCASCAN_N29_present_state_1_,
	FE_PT3_,
	FE_PT4_,
	SPCASCAN_N30_ov,
	SPCASCAN_N31_tdsp_state_2_,
	SPCASCAN_N32_two_cycle,
	SPCASCAN_N33_samp_int,
	n_7866,
	SPCASCAN_N35_three_cycle,
	dec_go_data,
	dec_go_prog,
	SPCASCAN_N36_tdsp_state_1_,
	n_7862);
   input SPCASCAN_N6_present_state_2_;
   input SPCASCAN_N7_present_state_1_;
   input FE_PT1_;
   input SPCASCAN_N23_done;
   input SPCASCAN_N28_read;
   input port_as;
   input FE_PT2_;
   input dec_go_port;
   input SPCASCAN_N29_present_state_1_;
   input FE_PT3_;
   input FE_PT4_;
   output SPCASCAN_N30_ov;
   input SPCASCAN_N31_tdsp_state_2_;
   output SPCASCAN_N32_two_cycle;
   input SPCASCAN_N33_samp_int;
   input n_7866;
   output SPCASCAN_N35_three_cycle;
   input dec_go_data;
   input dec_go_prog;
   input SPCASCAN_N36_tdsp_state_1_;
   input n_7862;

	input clk;
	input reset;
	input phi_1;
	input phi_2;
	input phi_3;
	input phi_4;
	input phi_5;
	input phi_6;
	input decode_skip_one;
	input gez;
	input gz;
	input nz;
	input z;
	input lz;
	input lez;
	output ov;
	input arnz;
	input bioz;
	input [32:0] alu_result;
	input [31:0] mpy_result;
	input [15:0] mdr;
	input [15:0] pdr;
	input [15:0] ir;
	input [15:0] decode;
	input [15:0] ar;
	output skip_one;
	output fetch_branch;
	output branch_stall;
	output pc_acc;
	output dmov_inc;
	output dp;
	output arp;
	output [15:0] ar0;
	output [15:0] ar1;
	output [15:0] pc;
	output [32:0] acc;
	output [31:0] p;
	output [15:0] top;
	output [3:0] alu_cmd;
	output [2:0] sel_op_a;
	output [2:0] sel_op_b;
	output read_prog;
	output go_prog;
	output read_data;
	output go_data;
	output read_port;
	output go_port;
	output ovm;
	input scan_en;
	input BG_scan_in;
	output BG_scan_out;

	wire [15:0] nbus_431;
	wire [2:0] nbus_435;
	wire [15:0] nbus_437;
	wire [2:0] nbus_439;



	INVXL i_10645(
		.A(n_7897),
		.Y(BG_scan_out));

	INVXL i_10644(
		.A(ar1[15]),
		.Y(n_7897));

	BUFX3 i_10360(
		.A(n_896),
		.Y(n_7516));

	CLKBUFX3 i_10358(
		.A(\nbus_436[0] ),
		.Y(n_7513));

	CLKBUFXL i_10357(
		.A(n_896),
		.Y(n_7510));

	CLKBUFXL i_10279(
		.A(\nbus_426[0] ),
		.Y(n_7423));

	CLKBUFXL i_10252(
		.A(\nbus_440[0] ),
		.Y(n_7384));

	CLKBUFXL i_10230(
		.A(\nbus_440[0] ),
		.Y(n_7353));

	BUFX2 i_10131(
		.A(n_794),
		.Y(n_7218));

	CLKBUFX2 i_10123(
		.A(n_1008),
		.Y(n_7206));

	CLKBUFX2 i_10121(
		.A(n_992),
		.Y(n_7203));

	CLKBUFX2 i_10119(
		.A(ir[12]),
		.Y(n_7200));

	BUFX3 i_10116(
		.A(n_7029),
		.Y(n_7197));

	CLKBUFXL i_10115(
		.A(n_1086),
		.Y(n_7194));

	CLKBUFXL i_10113(
		.A(n_1084),
		.Y(n_7191));

	CLKBUFXL i_10027(
		.A(ir[11]),
		.Y(n_7072));

	CLKBUFXL i_10007(
		.A(n_4221),
		.Y(n_7035));

	CLKBUFXL i_10004(
		.A(n_920),
		.Y(n_7029));

	CLKBUFXL i_10000(
		.A(\nbus_430[0] ),
		.Y(n_7021));

	CLKBUFXL i_9961(
		.A(\nbus_682[0] ),
		.Y(alu_cmd[0]));

	CLKBUFXL i_9957(
		.A(\nbus_681[1] ),
		.Y(alu_cmd[1]));

	CLKBUFXL i_9893(
		.A(\nbus_426[0] ),
		.Y(n_6812));

	CLKBUFXL i_9891(
		.A(\nbus_432[0] ),
		.Y(n_6809));

	CLKBUFX3 i_9525(
		.A(n_4221),
		.Y(n_6303));

	NAND2X1 i_579(
		.A(mdr[14]),
		.B(n_7029),
		.Y(n_600));

	NOR2X1 i_575(
		.A(ar[14]),
		.B(n_1031),
		.Y(n_595));

	OAI221XL i_248240(
		.A0(n_718),
		.A1(n_7206),
		.B0(n_720),
		.B1(n_7203),
		.C0(n_593),
		.Y(nbus_431[15]));

	NAND2X1 i_569(
		.A(mdr[15]),
		.B(n_7029),
		.Y(n_593));

	NOR2X1 i_567(
		.A(ar[15]),
		.B(n_1006),
		.Y(n_590));

	AOI32X1 i_2507(
		.A0(n_7218),
		.A1(n_850),
		.A2(n_792),
		.B0(n_855),
		.B1(n_4089),
		.Y(n_2082));

	NAND2X1 i_3501(
		.A(n_585),
		.B(n_474),
		.Y(\nbus_432[0] ));

	NAND3BX1 i_551(
		.AN(n_924),
		.B(n_809),
		.C(n_989),
		.Y(n_585));

	NAND2BX1 i_196(
		.AN(nbus_435[2]),
		.B(n_954),
		.Y(nbus_435[1]));

	NAND4BXL i_195(
		.AN(n_584),
		.B(n_934),
		.C(n_936),
		.D(n_926),
		.Y(nbus_435[2]));

	NOR3BX1 i_1694(
		.AN(ir[15]),
		.B(ir[13]),
		.C(ir[14]),
		.Y(n_584));

	AOI32X1 i_2445(
		.A0(ir[0]),
		.A1(n_893),
		.A2(n_871),
		.B0(mdr[0]),
		.B1(n_844),
		.Y(n_2534));

	AOI31X1 i_2440(
		.A0(n_7218),
		.A1(n_828),
		.A2(n_4090),
		.B0(n_399),
		.Y(n_2610));

	OAI21XL i_398239(
		.A0(n_7510),
		.A1(pc[0]),
		.B0(n_580),
		.Y(nbus_437[0]));

	NAND2X1 i_536(
		.A(decode[0]),
		.B(n_896),
		.Y(n_580));

	OAI21XL i_388238(
		.A0(n_7510),
		.A1(n_578),
		.B0(n_576),
		.Y(nbus_437[1]));

	XNOR2X1 i_244(
		.A(pc[1]),
		.B(pc[0]),
		.Y(n_578));

	NAND2X1 i_532(
		.A(decode[1]),
		.B(n_896),
		.Y(n_576));

	OAI21XL i_378237(
		.A0(n_7510),
		.A1(n_573),
		.B0(n_571),
		.Y(nbus_437[2]));

	AOI21X1 i_243(
		.A0(pc[2]),
		.A1(n_966),
		.B0(n_570),
		.Y(n_573));

	NAND2X1 i_527(
		.A(decode[2]),
		.B(n_896),
		.Y(n_571));

	NOR2X1 i_526(
		.A(pc[2]),
		.B(n_966),
		.Y(n_570));

	OAI21XL i_368236(
		.A0(n_7510),
		.A1(n_568),
		.B0(n_566),
		.Y(nbus_437[3]));

	AOI21X1 i_242(
		.A0(pc[3]),
		.A1(n_967),
		.B0(n_565),
		.Y(n_568));

	NAND2X1 i_522(
		.A(decode[3]),
		.B(n_896),
		.Y(n_566));

	NOR2X1 i_521(
		.A(pc[3]),
		.B(n_967),
		.Y(n_565));

	OAI21XL i_358235(
		.A0(n_896),
		.A1(n_563),
		.B0(n_561),
		.Y(nbus_437[4]));

	AOI21X1 i_241(
		.A0(pc[4]),
		.A1(n_968),
		.B0(n_560),
		.Y(n_563));

	NAND2X1 i_517(
		.A(decode[4]),
		.B(n_896),
		.Y(n_561));

	NOR2X1 i_516(
		.A(pc[4]),
		.B(n_968),
		.Y(n_560));

	OAI21XL i_348234(
		.A0(n_7510),
		.A1(n_558),
		.B0(n_556),
		.Y(nbus_437[5]));

	AOI21X1 i_240(
		.A0(pc[5]),
		.A1(n_969),
		.B0(n_555),
		.Y(n_558));

	NAND2X1 i_512(
		.A(decode[5]),
		.B(n_7516),
		.Y(n_556));

	NOR2X1 i_511(
		.A(pc[5]),
		.B(n_969),
		.Y(n_555));

	OAI21XL i_338233(
		.A0(n_7510),
		.A1(n_553),
		.B0(n_551),
		.Y(nbus_437[6]));

	AOI21X1 i_239(
		.A0(pc[6]),
		.A1(n_970),
		.B0(n_550),
		.Y(n_553));

	NAND2X1 i_507(
		.A(decode[6]),
		.B(n_7516),
		.Y(n_551));

	NOR2X1 i_506(
		.A(pc[6]),
		.B(n_970),
		.Y(n_550));

	OAI21XL i_32(
		.A0(n_7510),
		.A1(n_548),
		.B0(n_546),
		.Y(nbus_437[7]));

	AOI21X1 i_238(
		.A0(pc[7]),
		.A1(n_971),
		.B0(n_545),
		.Y(n_548));

	NAND2X1 i_502(
		.A(decode[7]),
		.B(n_7516),
		.Y(n_546));

	NOR2X1 i_501(
		.A(pc[7]),
		.B(n_971),
		.Y(n_545));

	OAI21XL i_318232(
		.A0(n_7510),
		.A1(n_543),
		.B0(n_541),
		.Y(nbus_437[8]));

	AOI21X1 i_237(
		.A0(pc[8]),
		.A1(n_972),
		.B0(n_540),
		.Y(n_543));

	NAND2X1 i_497(
		.A(decode[8]),
		.B(n_7516),
		.Y(n_541));

	NOR2X1 i_496(
		.A(pc[8]),
		.B(n_972),
		.Y(n_540));

	OAI21XL i_308231(
		.A0(n_7510),
		.A1(n_538),
		.B0(n_536),
		.Y(nbus_437[9]));

	AOI21X1 i_236(
		.A0(pc[9]),
		.A1(n_973),
		.B0(n_535),
		.Y(n_538));

	NAND2X1 i_492(
		.A(decode[9]),
		.B(n_7516),
		.Y(n_536));

	NOR2X1 i_491(
		.A(pc[9]),
		.B(n_973),
		.Y(n_535));

	OAI21XL i_298230(
		.A0(n_7510),
		.A1(n_533),
		.B0(n_531),
		.Y(nbus_437[10]));

	AOI21X1 i_235(
		.A0(pc[10]),
		.A1(n_974),
		.B0(n_529),
		.Y(n_533));

	NAND2X1 i_487(
		.A(decode[10]),
		.B(n_896),
		.Y(n_531));

	NOR2X1 i_485(
		.A(pc[10]),
		.B(n_974),
		.Y(n_529));

	OAI21XL i_288229(
		.A0(n_7510),
		.A1(n_528),
		.B0(n_526),
		.Y(nbus_437[11]));

	AOI21X1 i_234(
		.A0(pc[11]),
		.A1(n_975),
		.B0(n_524),
		.Y(n_528));

	NAND2X1 i_482(
		.A(decode[11]),
		.B(n_896),
		.Y(n_526));

	NOR2X1 i_480(
		.A(pc[11]),
		.B(n_975),
		.Y(n_524));

	MXI2X1 i_278228(
		.S0(n_7510),
		.B(decode[12]),
		.A(n_523),
		.Y(nbus_437[12]));

	OAI31X1 i_233(
		.A0(n_973),
		.A1(n_982),
		.A2(pc[12]),
		.B0(n_519),
		.Y(n_523));

	OAI21XL i_475(
		.A0(n_973),
		.A1(n_982),
		.B0(pc[12]),
		.Y(n_519));

	OAI21XL i_268227(
		.A0(n_7510),
		.A1(n_518),
		.B0(n_516),
		.Y(nbus_437[13]));

	XNOR2X1 i_232(
		.A(pc[13]),
		.B(n_984),
		.Y(n_518));

	NAND2X1 i_472(
		.A(decode[13]),
		.B(n_896),
		.Y(n_516));

	OAI21XL i_258226(
		.A0(n_7510),
		.A1(n_513),
		.B0(n_511),
		.Y(nbus_437[14]));

	XNOR2X1 i_231(
		.A(pc[14]),
		.B(n_981),
		.Y(n_513));

	NAND2X1 i_467(
		.A(decode[14]),
		.B(n_896),
		.Y(n_511));

	OAI21XL i_248225(
		.A0(n_508),
		.A1(n_7510),
		.B0(n_506),
		.Y(nbus_437[15]));

	XNOR2X1 i_230(
		.A(pc[15]),
		.B(n_978),
		.Y(n_508));

	NAND2X1 i_462(
		.A(decode[15]),
		.B(n_896),
		.Y(n_506));

	NAND2X1 i_2796(
		.A(phi_6),
		.B(SPCASCAN_N35_three_cycle),
		.Y(n_2768));

	OR4X1 i_1818651(
		.A(n_584),
		.B(n_871),
		.C(n_935),
		.D(n_496),
		.Y(nbus_439[0]));

	OAI21XL i_3732(
		.A0(n_503),
		.A1(n_959),
		.B0(\nbus_428[0] ),
		.Y(\nbus_434[0] ));

	AOI211X1 i_222(
		.A0(n_796),
		.A1(n_4082),
		.B0(n_952),
		.C0(n_584),
		.Y(n_503));

	AOI211X1 i_185(
		.A0(n_811),
		.A1(n_960),
		.B0(n_497),
		.C0(n_499),
		.Y(\nbus_428[0] ));

	AOI31X1 i_450(
		.A0(n_380),
		.A1(n_879),
		.A2(n_940),
		.B0(n_959),
		.Y(n_499));

	NOR3X1 i_446(
		.A(n_922),
		.B(n_829),
		.C(n_804),
		.Y(n_497));

	NAND4BXL i_1808650(
		.AN(n_955),
		.B(n_950),
		.C(n_936),
		.D(n_954),
		.Y(nbus_439[1]));

	AND3X1 i_441(
		.A(ir[15]),
		.B(ir[14]),
		.C(n_829),
		.Y(n_496));

	NAND2BX1 i_1798649(
		.AN(ir[15]),
		.B(n_494),
		.Y(nbus_439[2]));

	OAI31X1 i_438(
		.A0(n_952),
		.A1(n_820),
		.A2(n_951),
		.B0(ir[14]),
		.Y(n_494));

	AOI22X1 i_4078(
		.A0(n_948),
		.A1(n_949),
		.B0(n_941),
		.B1(n_491),
		.Y(n_2909));

	AOI21X1 i_179(
		.A0(ir[5]),
		.A1(ir[4]),
		.B0(n_478),
		.Y(n_493));

	NAND4X1 i_221(
		.A(n_945),
		.B(n_943),
		.C(n_489),
		.D(n_484),
		.Y(n_491));

	OAI21XL i_428(
		.A0(n_802),
		.A1(n_482),
		.B0(n_4080),
		.Y(n_489));

	OAI21XL i_178(
		.A0(ir[9]),
		.A1(n_788),
		.B0(n_481),
		.Y(n_485));

	NAND2X1 i_425(
		.A(n_871),
		.B(n_912),
		.Y(n_484));

	AOI211X1 i_124(
		.A0(ir[9]),
		.A1(ir[8]),
		.B0(ir[10]),
		.C0(n_913),
		.Y(n_483));

	NOR3X1 i_423(
		.A(n_889),
		.B(n_863),
		.C(n_483),
		.Y(n_482));

	NAND2X1 i_422(
		.A(n_7072),
		.B(n_800),
		.Y(n_481));

	NOR2X1 i_419(
		.A(ir[5]),
		.B(ir[4]),
		.Y(n_478));

	NAND2BX1 i_4136(
		.AN(n_475),
		.B(n_474),
		.Y(\nbus_440[0] ));

	AOI21X1 i_416(
		.A0(n_940),
		.A1(n_882),
		.B0(n_924),
		.Y(n_475));

	NAND2X1 i_415(
		.A(n_923),
		.B(n_811),
		.Y(n_474));

	NOR2X1 i_408(
		.A(n_863),
		.B(n_842),
		.Y(n_470));

	NOR2BX1 i_404(
		.AN(n_875),
		.B(n_868),
		.Y(n_467));

	AOI22X1 i_4206(
		.A0(n_466),
		.A1(n_4220),
		.B0(n_464),
		.B1(n_910),
		.Y(n_3146));

	NAND2BX1 i_218(
		.AN(n_7197),
		.B(n_462),
		.Y(n_466));

	NAND4X1 i_219(
		.A(n_917),
		.B(n_461),
		.C(n_456),
		.D(n_912),
		.Y(n_464));

	NAND3BX1 i_399(
		.AN(update_stall),
		.B(phi_6),
		.C(n_1105),
		.Y(n_462));

	NAND2X1 i_389(
		.A(SPCASCAN_N35_three_cycle),
		.B(n_828),
		.Y(n_461));

	OAI21XL i_392(
		.A0(n_813),
		.A1(SPCASCAN_N32_two_cycle),
		.B0(n_809),
		.Y(n_456));

	OAI221XL i_227(
		.A0(n_7072),
		.A1(ir[10]),
		.B0(n_791),
		.B1(n_788),
		.C0(n_800),
		.Y(n_455));

	NAND3X1 i_380(
		.A(n_908),
		.B(n_877),
		.C(n_875),
		.Y(n_450));

	OAI221XL i_3965(
		.A0(n_448),
		.A1(n_905),
		.B0(n_831),
		.B1(n_814),
		.C0(n_404),
		.Y(n_2765));

	AOI21X1 i_183(
		.A0(n_446),
		.A1(n_4092),
		.B0(n_828),
		.Y(n_448));

	OAI21XL i_79(
		.A0(n_804),
		.A1(n_829),
		.B0(n_401),
		.Y(n_447));

	NAND2X1 i_133(
		.A(n_813),
		.B(n_804),
		.Y(n_446));

	OAI21XL i_3880(
		.A0(n_444),
		.A1(n_797),
		.B0(n_896),
		.Y(\nbus_436[0] ));

	AOI221X1 i_35(
		.A0(SPCASCAN_N30_ov),
		.A1(n_839),
		.B0(n_440),
		.B1(n_836),
		.C0(n_442),
		.Y(n_444));

	NOR2BX1 i_367(
		.AN(n_835),
		.B(n_438),
		.Y(n_442));

	OAI2BB1X1 i_248(
		.A0N(bioz),
		.A1N(n_791),
		.B0(n_899),
		.Y(n_440));

	AOI211X1 i_249(
		.A0(gez),
		.A1(n_4084),
		.B0(n_902),
		.C0(n_430),
		.Y(n_438));

	NAND3X1 i_353(
		.A(n_841),
		.B(n_4085),
		.C(lz),
		.Y(n_432));

	NAND3X1 i_354(
		.A(lez),
		.B(n_843),
		.C(n_4085),
		.Y(n_431));

	NOR2BX1 i_351(
		.AN(n_844),
		.B(nz),
		.Y(n_430));

	OR2X1 i_180(
		.A(n_893),
		.B(n_844),
		.Y(n_429));

	AOI21X1 i_3737(
		.A0(phi_6),
		.A1(branch_stall_delay),
		.B0(n_4083),
		.Y(n_2515));

	AOI211X1 i_3576(
		.A0(alu_result[32]),
		.A1(n_425),
		.B0(n_427),
		.C0(n_423),
		.Y(n_2384));

	AND4X1 i_343(
		.A(phi_1),
		.B(n_7218),
		.C(SPCASCAN_N30_ov),
		.D(n_839),
		.Y(n_427));

	OAI2BB2X1 i_212(
		.A0N(n_811),
		.A1N(n_4089),
		.B0(n_805),
		.B1(n_890),
		.Y(n_425));

	NAND4BXL i_213(
		.AN(n_823),
		.B(n_886),
		.C(n_883),
		.D(n_882),
		.Y(n_424));

	AND4X1 i_341(
		.A(phi_6),
		.B(n_7218),
		.C(alu_result[32]),
		.D(n_424),
		.Y(n_423));

	NOR2X1 i_3659(
		.A(n_1106),
		.B(phi_3),
		.Y(n_2115));

	AOI2BB1X1 i_3351(
		.A0N(n_414),
		.A1N(n_830),
		.B0(phi_3),
		.Y(n_2079));

	AOI21X1 i_210(
		.A0(n_787),
		.A1(n_792),
		.B0(n_855),
		.Y(n_414));

	NOR4BX1 i_3842(
		.AN(n_410),
		.B(n_409),
		.C(phi_3),
		.D(n_399),
		.Y(n_1940));

	NAND2BX1 i_305(
		.AN(n_784),
		.B(n_395),
		.Y(n_410));

	NOR2X1 i_302(
		.A(n_790),
		.B(n_851),
		.Y(n_409));

	OAI211X1 i_295(
		.A0(n_383),
		.A1(phi_1),
		.B0(n_7218),
		.C0(n_835),
		.Y(n_407));

	NAND2X1 i_290(
		.A(n_4085),
		.B(n_835),
		.Y(n_406));

	NOR4BX1 i_3157(
		.AN(n_404),
		.B(n_405),
		.C(n_403),
		.D(n_2235),
		.Y(n_1833));

	NOR2X1 i_285(
		.A(n_804),
		.B(n_830),
		.Y(n_405));

	NAND2X1 i_284(
		.A(n_7218),
		.B(n_447),
		.Y(n_404));

	AOI21X1 i_283(
		.A0(n_816),
		.A1(n_793),
		.B0(n_830),
		.Y(n_403));

	NAND2X1 i_280(
		.A(n_828),
		.B(n_4090),
		.Y(n_401));

	OR2X1 i_3483(
		.A(n_400),
		.B(n_399),
		.Y(n_2235));

	NOR2X1 i_275(
		.A(n_814),
		.B(n_831),
		.Y(n_400));

	NOR2X1 i_274(
		.A(n_813),
		.B(n_830),
		.Y(n_399));

	AOI222X1 i_3117(
		.A0(skip_one),
		.A1(phi_1),
		.B0(n_396),
		.B1(n_395),
		.C0(n_796),
		.C1(n_697),
		.Y(n_1790));

	NAND3BX1 i_209(
		.AN(n_817),
		.B(n_818),
		.C(n_699),
		.Y(n_396));

	AOI211X1 i_52(
		.A0(n_793),
		.A1(n_816),
		.B0(branch_stall_delay),
		.C0(branch_stall),
		.Y(n_395));

	NAND2BX1 i_2462(
		.AN(n_584),
		.B(n_2387),
		.Y(nbus_435[0]));

	AOI211X1 i_2797(
		.A0(ir[14]),
		.A1(n_4078),
		.B0(n_807),
		.C0(n_802),
		.Y(n_2387));

	OAI32X1 i_2874(
		.A0(n_797),
		.A1(n_793),
		.A2(n_4077),
		.B0(n_784),
		.B1(n_795),
		.Y(n_1439));

	NOR3BX1 i_1731(
		.AN(n_847),
		.B(n_839),
		.C(n_836),
		.Y(n_383));

	NAND2BX1 i_63(
		.AN(n_913),
		.B(n_4079),
		.Y(n_382));

	NAND3X1 i_2232(
		.A(ir[2]),
		.B(ir[0]),
		.C(n_869),
		.Y(n_380));

	OAI221XL i_258241(
		.A0(n_722),
		.A1(n_7206),
		.B0(n_724),
		.B1(n_7203),
		.C0(n_600),
		.Y(nbus_431[14]));

	NOR2X1 i_586(
		.A(ar[13]),
		.B(n_1036),
		.Y(n_602));

	NAND2X1 i_589(
		.A(mdr[13]),
		.B(n_7029),
		.Y(n_606));

	OAI221XL i_268242(
		.A0(n_726),
		.A1(n_7206),
		.B0(n_728),
		.B1(n_7203),
		.C0(n_606),
		.Y(nbus_431[13]));

	NAND2X1 i_597(
		.A(mdr[12]),
		.B(n_7029),
		.Y(n_612));

	OAI221XL i_278243(
		.A0(n_730),
		.A1(n_7206),
		.B0(n_732),
		.B1(n_7203),
		.C0(n_612),
		.Y(nbus_431[12]));

	NOR2X1 i_602(
		.A(ar[11]),
		.B(n_1018),
		.Y(n_614));

	NAND2X1 i_606(
		.A(mdr[11]),
		.B(n_7197),
		.Y(n_619));

	OAI221XL i_288244(
		.A0(n_734),
		.A1(n_7206),
		.B0(n_736),
		.B1(n_7203),
		.C0(n_619),
		.Y(nbus_431[11]));

	NOR2X1 i_611(
		.A(ar[10]),
		.B(n_1017),
		.Y(n_621));

	NAND2X1 i_614(
		.A(mdr[10]),
		.B(n_7029),
		.Y(n_625));

	OAI221XL i_298245(
		.A0(n_738),
		.A1(n_7206),
		.B0(n_740),
		.B1(n_7203),
		.C0(n_625),
		.Y(nbus_431[10]));

	NOR2X1 i_619(
		.A(ar[9]),
		.B(n_1033),
		.Y(n_627));

	NAND2X1 i_622(
		.A(mdr[9]),
		.B(n_7197),
		.Y(n_631));

	OAI221XL i_308246(
		.A0(n_742),
		.A1(n_7206),
		.B0(n_744),
		.B1(n_7203),
		.C0(n_631),
		.Y(nbus_431[9]));

	OAI21XL i_627(
		.A0(n_4073),
		.A1(ar[7]),
		.B0(ar[8]),
		.Y(n_633));

	NOR2X1 i_629(
		.A(ar[8]),
		.B(n_1015),
		.Y(n_635));

	NAND2X1 i_630(
		.A(mdr[8]),
		.B(n_7197),
		.Y(n_637));

	OAI221XL i_318247(
		.A0(n_748),
		.A1(n_7206),
		.B0(n_747),
		.B1(n_7203),
		.C0(n_637),
		.Y(nbus_431[8]));

	NOR2X1 i_636(
		.A(ar[7]),
		.B(n_1014),
		.Y(n_640));

	NOR2X1 i_640(
		.A(n_750),
		.B(n_7206),
		.Y(n_644));

	NAND2X1 i_328248(
		.A(n_1044),
		.B(n_1045),
		.Y(nbus_431[7]));

	NOR2X1 i_645(
		.A(ar[6]),
		.B(n_1013),
		.Y(n_647));

	NOR2X1 i_649(
		.A(n_754),
		.B(n_7206),
		.Y(n_651));

	NAND2X1 i_338249(
		.A(n_1046),
		.B(n_1047),
		.Y(nbus_431[6]));

	OAI21XL i_653(
		.A0(n_4074),
		.A1(ar[4]),
		.B0(ar[5]),
		.Y(n_653));

	NOR2X1 i_655(
		.A(ar[5]),
		.B(n_1012),
		.Y(n_655));

	NOR2X1 i_658(
		.A(n_758),
		.B(n_7203),
		.Y(n_658));

	NAND2X1 i_348250(
		.A(n_1048),
		.B(n_1049),
		.Y(nbus_431[5]));

	NOR2X1 i_662(
		.A(ar[4]),
		.B(n_1011),
		.Y(n_660));

	NOR2X1 i_667(
		.A(n_762),
		.B(n_7206),
		.Y(n_665));

	NAND2X1 i_358251(
		.A(n_1050),
		.B(n_1051),
		.Y(nbus_431[4]));

	NOR2X1 i_672(
		.A(ar[3]),
		.B(n_1010),
		.Y(n_668));

	NOR2X1 i_676(
		.A(n_766),
		.B(n_7206),
		.Y(n_672));

	NAND2X1 i_368252(
		.A(n_1052),
		.B(n_1053),
		.Y(nbus_431[3]));

	NOR2X1 i_681(
		.A(n_1009),
		.B(ar[2]),
		.Y(n_675));

	OAI21XL i_682(
		.A0(ar[0]),
		.A1(ar[1]),
		.B0(ar[2]),
		.Y(n_676));

	NOR2X1 i_685(
		.A(n_770),
		.B(n_7206),
		.Y(n_679));

	NAND2X1 i_378253(
		.A(n_1054),
		.B(n_1055),
		.Y(nbus_431[2]));

	NAND2X1 i_388254(
		.A(n_1056),
		.B(n_1058),
		.Y(nbus_431[1]));

	NAND4X1 i_696(
		.A(n_7072),
		.B(n_7200),
		.C(n_821),
		.D(n_4079),
		.Y(n_686));

	NAND2BX1 i_699(
		.AN(n_693),
		.B(n_948),
		.Y(n_687));

	OAI21XL i_223(
		.A0(n_863),
		.A1(n_4080),
		.B0(n_686),
		.Y(n_689));

	OAI2BB1X1 i_3282(
		.A0N(n_689),
		.A1N(n_941),
		.B0(n_687),
		.Y(\nbus_430[0] ));

	AND2X1 i_136(
		.A(n_1008),
		.B(n_992),
		.Y(n_693));

	OAI21XL i_398255(
		.A0(n_693),
		.A1(ar[0]),
		.B0(n_1061),
		.Y(nbus_431[0]));

	NOR2BX1 i_2655(
		.AN(n_2610),
		.B(n_409),
		.Y(n_1943));

	OAI22X1 i_76(
		.A0(n_814),
		.A1(n_4220),
		.B0(n_804),
		.B1(n_805),
		.Y(n_697));

	NAND2X1 i_55(
		.A(phi_4),
		.B(SPCASCAN_N35_three_cycle),
		.Y(n_699));

	AOI22X1 i_228(
		.A0(n_816),
		.A1(n_793),
		.B0(n_1064),
		.B1(n_830),
		.Y(n_700));

	AOI22X1 i_2385(
		.A0(n_700),
		.A1(n_699),
		.B0(n_697),
		.B1(n_796),
		.Y(n_1793));

	OR3XL i_1798667(
		.A(n_925),
		.B(n_937),
		.C(n_1065),
		.Y(\nbus_429[2] ));

	NOR4BX1 i_1808668(
		.AN(n_926),
		.B(n_821),
		.C(n_937),
		.D(n_932),
		.Y(\nbus_429[1] ));

	NAND2X1 i_722(
		.A(n_809),
		.B(n_884),
		.Y(n_701));

	NOR3X1 i_203(
		.A(ir[10]),
		.B(n_4100),
		.C(n_872),
		.Y(n_704));

	AOI21X1 i_726(
		.A0(n_872),
		.A1(n_701),
		.B0(n_806),
		.Y(n_705));

	OAI32X1 i_2924(
		.A0(n_922),
		.A1(n_818),
		.A2(n_804),
		.B0(n_924),
		.B1(n_962),
		.Y(\nbus_426[0] ));

	AOI21X1 i_73(
		.A0(n_788),
		.A1(n_806),
		.B0(n_840),
		.Y(n_710));

	NOR2X1 i_747(
		.A(n_931),
		.B(n_1076),
		.Y(n_712));

	OAI32X1 i_112(
		.A0(n_841),
		.A1(n_844),
		.A2(n_4087),
		.B0(n_710),
		.B1(n_4086),
		.Y(n_713));

	OAI21XL i_743(
		.A0(n_821),
		.A1(n_808),
		.B0(n_7200),
		.Y(n_714));

	NAND2X1 i_744(
		.A(n_802),
		.B(n_4080),
		.Y(n_715));

	NAND3BX1 i_745(
		.AN(n_989),
		.B(n_809),
		.C(n_813),
		.Y(n_716));

	NOR3X1 i_746(
		.A(n_935),
		.B(n_951),
		.C(n_863),
		.Y(n_717));

	XNOR2X1 i_83(
		.A(ar[15]),
		.B(n_1022),
		.Y(n_718));

	AOI21X1 i_84(
		.A0(ar[15]),
		.A1(n_1006),
		.B0(n_590),
		.Y(n_720));

	OAI221XL i_248256(
		.A0(n_7194),
		.A1(n_718),
		.B0(n_7191),
		.B1(n_720),
		.C0(n_593),
		.Y(\nbus_425[15] ));

	AOI21X1 i_85(
		.A0(ar[14]),
		.A1(n_1031),
		.B0(n_595),
		.Y(n_722));

	XNOR2X1 i_86(
		.A(ar[14]),
		.B(n_1027),
		.Y(n_724));

	OAI221XL i_258257(
		.A0(n_7194),
		.A1(n_722),
		.B0(n_7191),
		.B1(n_724),
		.C0(n_600),
		.Y(\nbus_425[14] ));

	AOI21X1 i_87(
		.A0(ar[13]),
		.A1(n_1036),
		.B0(n_602),
		.Y(n_726));

	AOI21X1 i_88(
		.A0(ar[13]),
		.A1(n_4075),
		.B0(n_1027),
		.Y(n_728));

	OAI221XL i_268258(
		.A0(n_7194),
		.A1(n_726),
		.B0(n_728),
		.B1(n_7191),
		.C0(n_606),
		.Y(\nbus_425[13] ));

	XNOR2X1 i_89(
		.A(ar[12]),
		.B(n_1029),
		.Y(n_730));

	AOI21X1 i_90(
		.A0(ar[12]),
		.A1(n_1025),
		.B0(n_1026),
		.Y(n_732));

	OAI221XL i_278259(
		.A0(n_7194),
		.A1(n_730),
		.B0(n_7191),
		.B1(n_732),
		.C0(n_612),
		.Y(\nbus_425[12] ));

	AOI21X1 i_91(
		.A0(ar[11]),
		.A1(n_1018),
		.B0(n_614),
		.Y(n_734));

	XNOR2X1 i_92(
		.A(ar[11]),
		.B(n_1002),
		.Y(n_736));

	OAI221XL i_288260(
		.A0(n_7194),
		.A1(n_734),
		.B0(n_7191),
		.B1(n_736),
		.C0(n_619),
		.Y(\nbus_425[11] ));

	AOI21X1 i_93(
		.A0(ar[10]),
		.A1(n_1017),
		.B0(n_621),
		.Y(n_738));

	AOI21X1 i_94(
		.A0(ar[10]),
		.A1(n_4072),
		.B0(n_1002),
		.Y(n_740));

	OAI221XL i_298261(
		.A0(n_7194),
		.A1(n_738),
		.B0(n_740),
		.B1(n_7191),
		.C0(n_625),
		.Y(\nbus_425[10] ));

	AOI21X1 i_95(
		.A0(ar[9]),
		.A1(n_1033),
		.B0(n_627),
		.Y(n_742));

	AOI21X1 i_96(
		.A0(ar[9]),
		.A1(n_1000),
		.B0(n_1001),
		.Y(n_744));

	OAI221XL i_308262(
		.A0(n_7194),
		.A1(n_742),
		.B0(n_7191),
		.B1(n_744),
		.C0(n_631),
		.Y(\nbus_425[9] ));

	AND2X1 i_97(
		.A(n_1000),
		.B(n_633),
		.Y(n_747));

	AOI21X1 i_106(
		.A0(ar[8]),
		.A1(n_1015),
		.B0(n_635),
		.Y(n_748));

	OAI221XL i_318263(
		.A0(n_7194),
		.A1(n_748),
		.B0(n_747),
		.B1(n_7191),
		.C0(n_637),
		.Y(\nbus_425[8] ));

	AOI21X1 i_99(
		.A0(ar[7]),
		.A1(n_1014),
		.B0(n_640),
		.Y(n_750));

	AOI21X1 i_100(
		.A0(ar[7]),
		.A1(n_4073),
		.B0(n_999),
		.Y(n_751));

	OAI221XL i_328264(
		.A0(n_751),
		.A1(n_7191),
		.B0(n_7194),
		.B1(n_750),
		.C0(n_1044),
		.Y(\nbus_425[7] ));

	AOI21X1 i_101(
		.A0(ar[6]),
		.A1(n_1013),
		.B0(n_647),
		.Y(n_754));

	AOI21X1 i_120(
		.A0(ar[6]),
		.A1(n_997),
		.B0(n_998),
		.Y(n_755));

	OAI221XL i_338265(
		.A0(n_7191),
		.A1(n_755),
		.B0(n_7194),
		.B1(n_754),
		.C0(n_1046),
		.Y(\nbus_425[6] ));

	AND2X1 i_102(
		.A(n_997),
		.B(n_653),
		.Y(n_758));

	AOI21X1 i_109(
		.A0(ar[5]),
		.A1(n_1012),
		.B0(n_655),
		.Y(n_759));

	OAI221XL i_348266(
		.A0(n_7194),
		.A1(n_759),
		.B0(n_758),
		.B1(n_7191),
		.C0(n_1048),
		.Y(\nbus_425[5] ));

	AOI21X1 i_103(
		.A0(ar[4]),
		.A1(n_1011),
		.B0(n_660),
		.Y(n_762));

	AOI21X1 i_121(
		.A0(ar[4]),
		.A1(n_4074),
		.B0(n_996),
		.Y(n_763));

	OAI221XL i_358267(
		.A0(n_763),
		.A1(n_7191),
		.B0(n_7194),
		.B1(n_762),
		.C0(n_1050),
		.Y(\nbus_425[4] ));

	AOI21X1 i_110(
		.A0(ar[3]),
		.A1(n_1010),
		.B0(n_668),
		.Y(n_766));

	AOI21X1 i_125(
		.A0(ar[3]),
		.A1(n_994),
		.B0(n_995),
		.Y(n_767));

	OAI221XL i_368268(
		.A0(n_7191),
		.A1(n_767),
		.B0(n_7194),
		.B1(n_766),
		.C0(n_1052),
		.Y(\nbus_425[3] ));

	AOI21X1 i_104(
		.A0(ar[2]),
		.A1(n_1009),
		.B0(n_675),
		.Y(n_770));

	AND2X1 i_122(
		.A(n_994),
		.B(n_676),
		.Y(n_771));

	OAI221XL i_378269(
		.A0(n_771),
		.A1(n_7191),
		.B0(n_7194),
		.B1(n_770),
		.C0(n_1054),
		.Y(\nbus_425[2] ));

	NAND2BX1 i_824(
		.AN(n_7191),
		.B(n_1057),
		.Y(n_774));

	OAI211X1 i_388270(
		.A0(n_7194),
		.A1(n_1057),
		.B0(n_1056),
		.C0(n_774),
		.Y(\nbus_425[1] ));

	NAND4BXL i_829(
		.AN(n_837),
		.B(n_7072),
		.C(n_7200),
		.D(n_821),
		.Y(n_777));

	OAI31X1 i_225(
		.A0(n_7072),
		.A1(n_837),
		.A2(n_863),
		.B0(n_777),
		.Y(n_780));

	AOI22X1 i_2811(
		.A0(n_780),
		.A1(n_941),
		.B0(n_782),
		.B1(n_948),
		.Y(\nbus_424[0] ));

	NAND2BX1 i_834(
		.AN(ar[0]),
		.B(n_782),
		.Y(n_781));

	NAND2X1 i_137(
		.A(n_1086),
		.B(n_1084),
		.Y(n_782));

	NOR2X1 i_71(
		.A(SPCASCAN_N35_three_cycle),
		.B(n_4092),
		.Y(n_783));

	NAND2X1 i_21022(
		.A(phi_6),
		.B(n_783),
		.Y(n_784));

	NAND2X1 i_38(
		.A(ir[15]),
		.B(ir[14]),
		.Y(n_785));

	NAND3X1 i_78(
		.A(ir[15]),
		.B(ir[14]),
		.C(ir[13]),
		.Y(n_786));

	NOR2X1 i_1701(
		.A(n_7200),
		.B(n_786),
		.Y(n_787));

	NAND2X1 i_23(
		.A(ir[10]),
		.B(ir[8]),
		.Y(n_788));

	NOR2X1 i_28(
		.A(ir[9]),
		.B(n_788),
		.Y(n_789));

	NAND2X1 i_115(
		.A(n_7072),
		.B(n_789),
		.Y(n_790));

	NOR2BX1 i_20(
		.AN(ir[9]),
		.B(n_7072),
		.Y(n_791));

	NOR2BX1 i_193(
		.AN(n_791),
		.B(n_788),
		.Y(n_792));

	OAI21XL i_0(
		.A0(n_792),
		.A1(n_4084),
		.B0(n_787),
		.Y(n_793));

	NOR2X1 i_29(
		.A(branch_stall_delay),
		.B(branch_stall),
		.Y(n_794));

	NAND2BX1 i_189(
		.AN(n_793),
		.B(n_7218),
		.Y(n_795));

	NOR2X1 i_44(
		.A(SPCASCAN_N35_three_cycle),
		.B(SPCASCAN_N32_two_cycle),
		.Y(n_796));

	NAND2X1 i_170(
		.A(n_7218),
		.B(phi_1),
		.Y(n_797));

	NOR2X1 i_62(
		.A(ir[10]),
		.B(ir[9]),
		.Y(n_799));

	NAND2X1 i_21(
		.A(n_799),
		.B(n_4100),
		.Y(n_800));

	NOR2X1 i_37(
		.A(n_7072),
		.B(n_800),
		.Y(n_801));

	NOR2X1 i_1765(
		.A(ir[13]),
		.B(n_785),
		.Y(n_802));

	NAND3BX1 i_22(
		.AN(n_7200),
		.B(n_802),
		.C(n_801),
		.Y(n_804));

	NAND2X1 i_67(
		.A(phi_3),
		.B(n_7218),
		.Y(n_805));

	NAND2X1 i_24(
		.A(ir[10]),
		.B(n_4100),
		.Y(n_806));

	NOR2X1 i_256(
		.A(ir[15]),
		.B(ir[13]),
		.Y(n_807));

	AND2X1 i_1756(
		.A(ir[14]),
		.B(n_807),
		.Y(n_808));

	NOR2BX1 i_1790(
		.AN(n_808),
		.B(n_7200),
		.Y(n_809));

	AND2X1 i_194(
		.A(n_809),
		.B(n_791),
		.Y(n_810));

	AND2X1 i_1845(
		.A(n_810),
		.B(n_4087),
		.Y(n_811));

	NOR3X1 i_45(
		.A(ir[9]),
		.B(n_788),
		.C(n_7072),
		.Y(n_812));

	AOI21X1 i_1808(
		.A0(n_809),
		.A1(n_812),
		.B0(n_811),
		.Y(n_813));

	NAND2BX1 i_200(
		.AN(n_813),
		.B(n_7218),
		.Y(n_814));

	NAND3BX1 i_1763(
		.AN(ir[14]),
		.B(ir[15]),
		.C(ir[13]),
		.Y(n_816));

	AOI21X1 i_27(
		.A0(SPCASCAN_N32_two_cycle),
		.A1(SPCASCAN_N35_three_cycle),
		.B0(n_4220),
		.Y(n_817));

	NAND2X1 i_21039(
		.A(phi_6),
		.B(n_796),
		.Y(n_818));

	NAND2BX1 i_11(
		.AN(ir[15]),
		.B(ir[13]),
		.Y(n_820));

	NOR2X1 i_1753(
		.A(ir[14]),
		.B(n_820),
		.Y(n_821));

	NOR3X1 i_1750(
		.A(ir[15]),
		.B(ir[13]),
		.C(ir[14]),
		.Y(n_823));

	NAND2X1 i_128(
		.A(ir[14]),
		.B(n_4078),
		.Y(n_824));

	NAND2X1 i_3(
		.A(n_793),
		.B(n_816),
		.Y(n_828));

	NAND2X1 i_21014(
		.A(phi_3),
		.B(n_783),
		.Y(n_829));

	NAND3X1 i_174(
		.A(phi_6),
		.B(n_7218),
		.C(n_796),
		.Y(n_830));

	NAND2X1 i_153(
		.A(phi_5),
		.B(n_783),
		.Y(n_831));

	NAND2X1 i_282(
		.A(n_7200),
		.B(n_4088),
		.Y(n_832));

	NOR2BX1 i_1702(
		.AN(n_7200),
		.B(n_786),
		.Y(n_835));

	AND2X1 i_77(
		.A(n_835),
		.B(n_4087),
		.Y(n_836));

	NAND2X1 i_31(
		.A(n_799),
		.B(ir[8]),
		.Y(n_837));

	NOR2BX1 i_172(
		.AN(n_7072),
		.B(n_837),
		.Y(n_838));

	AND2X1 i_207(
		.A(n_835),
		.B(n_838),
		.Y(n_839));

	NAND2X1 i_26(
		.A(ir[9]),
		.B(n_7072),
		.Y(n_840));

	NOR2X1 i_33(
		.A(ir[10]),
		.B(ir[8]),
		.Y(n_841));

	NAND2X1 i_171(
		.A(n_841),
		.B(n_4085),
		.Y(n_842));

	NOR2X1 i_43(
		.A(ir[10]),
		.B(n_4100),
		.Y(n_843));

	NOR2X1 i_50(
		.A(n_788),
		.B(n_840),
		.Y(n_844));

	NOR4BX1 i_293(
		.AN(n_406),
		.B(n_812),
		.C(n_844),
		.D(n_4084),
		.Y(n_847));

	NOR3X1 i_186(
		.A(n_7200),
		.B(n_786),
		.C(n_818),
		.Y(n_850));

	NAND2X1 i_188(
		.A(n_7218),
		.B(n_850),
		.Y(n_851));

	OAI21XL i_80(
		.A0(n_7200),
		.A1(n_816),
		.B0(n_813),
		.Y(n_855));

	NOR2BX1 i_318(
		.AN(update_it),
		.B(update_stall),
		.Y(n_856));

	NAND4X1 i_39(
		.A(ir[7]),
		.B(phi_6),
		.C(n_856),
		.D(n_4220),
		.Y(n_859));

	NAND3X1 i_1937(
		.A(ir[14]),
		.B(ir[12]),
		.C(n_4078),
		.Y(n_863));

	NAND2BX1 i_2207(
		.AN(n_863),
		.B(n_844),
		.Y(n_864));

	NOR2BX1 i_187(
		.AN(ir[7]),
		.B(ir[6]),
		.Y(n_865));

	NAND4BXL i_40(
		.AN(n_864),
		.B(ir[3]),
		.C(n_478),
		.D(n_865),
		.Y(n_868));

	NOR2BX1 i_206(
		.AN(ir[1]),
		.B(n_868),
		.Y(n_869));

	NOR2X1 i_1935(
		.A(n_824),
		.B(ir[12]),
		.Y(n_871));

	NAND2X1 i_41(
		.A(n_871),
		.B(n_791),
		.Y(n_872));

	NOR2X1 i_127(
		.A(ir[0]),
		.B(n_864),
		.Y(n_873));

	NOR4X1 i_162(
		.A(ir[0]),
		.B(n_864),
		.C(ir[1]),
		.D(ir[2]),
		.Y(n_875));

	NOR2BX1 i_205(
		.AN(ir[4]),
		.B(ir[5]),
		.Y(n_876));

	NOR2BX1 i_333(
		.AN(n_865),
		.B(ir[3]),
		.Y(n_877));

	AOI33X1 i_7(
		.A0(n_876),
		.A1(n_877),
		.A2(n_875),
		.B0(n_871),
		.B1(n_841),
		.B2(n_791),
		.Y(n_879));

	NAND2X1 i_60(
		.A(n_380),
		.B(n_879),
		.Y(n_880));

	AOI31X1 i_75(
		.A0(SPCASCAN_N35_three_cycle),
		.A1(n_4092),
		.A2(n_4082),
		.B0(n_880),
		.Y(n_882));

	AOI21X1 i_17(
		.A0(n_871),
		.A1(n_801),
		.B0(n_704),
		.Y(n_883));

	NOR2X1 i_160(
		.A(n_7072),
		.B(ir[9]),
		.Y(n_884));

	AOI32X1 i_8(
		.A0(n_884),
		.A1(n_809),
		.A2(n_4087),
		.B0(n_841),
		.B1(n_810),
		.Y(n_886));

	NOR2X1 i_47(
		.A(n_7072),
		.B(n_837),
		.Y(n_889));

	NAND2X1 i_2132(
		.A(n_889),
		.B(n_871),
		.Y(n_890));

	NOR2X1 i_201(
		.A(n_840),
		.B(n_806),
		.Y(n_893));

	NOR2X1 i_350(
		.A(SPCASCAN_N32_two_cycle),
		.B(skip_one),
		.Y(n_895));

	NAND2X1 i_21079(
		.A(phi_6),
		.B(n_895),
		.Y(n_896));

	NOR2BX1 i_363(
		.AN(gz),
		.B(ir[9]),
		.Y(n_897));

	AOI222X1 i_365(
		.A0(n_7072),
		.A1(n_897),
		.B0(arnz),
		.B1(n_884),
		.C0(nz),
		.C1(n_4085),
		.Y(n_899));

	NAND3BX1 i_357(
		.AN(n_812),
		.B(n_431),
		.C(n_432),
		.Y(n_902));

	NAND3X1 i_376(
		.A(phi_6),
		.B(n_7218),
		.C(SPCASCAN_N35_three_cycle),
		.Y(n_905));

	NOR2BX1 i_204(
		.AN(ir[5]),
		.B(ir[4]),
		.Y(n_908));

	NOR2X1 i_46(
		.A(n_1105),
		.B(phi_1),
		.Y(n_910));

	AOI22X1 i_1987(
		.A0(n_455),
		.A1(n_871),
		.B0(n_4086),
		.B1(n_4100),
		.Y(n_912));

	NAND2BX1 i_36(
		.AN(n_863),
		.B(n_7072),
		.Y(n_913));

	AOI21X1 i_393(
		.A0(n_7200),
		.A1(n_808),
		.B0(n_823),
		.Y(n_914));

	OAI21XL i_394(
		.A0(n_4092),
		.A1(n_804),
		.B0(n_914),
		.Y(n_915));

	AOI211X1 i_396(
		.A0(n_884),
		.A1(n_836),
		.B0(n_915),
		.C0(n_483),
		.Y(n_917));

	NOR3X1 i_6(
		.A(ir[14]),
		.B(n_1105),
		.C(n_820),
		.Y(n_920));

	NAND2X1 i_4(
		.A(n_794),
		.B(n_6303),
		.Y(n_922));

	NOR2X1 i_192(
		.A(n_922),
		.B(n_818),
		.Y(n_923));

	NAND2X1 i_51(
		.A(phi_6),
		.B(n_4076),
		.Y(n_924));

	NAND2BX1 i_18(
		.AN(n_467),
		.B(n_382),
		.Y(n_925));

	NAND2X1 i_1858(
		.A(n_843),
		.B(n_810),
		.Y(n_926));

	NAND2X1 i_118(
		.A(n_926),
		.B(n_886),
		.Y(n_927));

	AOI211X1 i_406(
		.A0(ir[13]),
		.A1(n_7200),
		.B0(ir[15]),
		.C0(ir[14]),
		.Y(n_928));

	NOR3X1 i_81(
		.A(n_927),
		.B(n_928),
		.C(n_925),
		.Y(n_930));

	NAND2X1 i_61(
		.A(n_890),
		.B(n_883),
		.Y(n_931));

	OAI21XL i_9(
		.A0(n_837),
		.A1(n_913),
		.B0(n_4091),
		.Y(n_932));

	AOI32X1 i_72(
		.A0(ir[2]),
		.A1(n_873),
		.A2(n_869),
		.B0(n_871),
		.B1(n_812),
		.Y(n_934));

	NOR2BX1 i_2194(
		.AN(n_893),
		.B(n_863),
		.Y(n_935));

	AOI21X1 i_119(
		.A0(n_4086),
		.A1(n_4087),
		.B0(n_935),
		.Y(n_936));

	NAND2X1 i_19(
		.A(n_934),
		.B(n_936),
		.Y(n_937));

	NOR4BX1 i_113(
		.AN(n_930),
		.B(n_937),
		.C(n_932),
		.D(n_931),
		.Y(n_940));

	NOR3X1 i_49(
		.A(n_1105),
		.B(phi_1),
		.C(reset),
		.Y(n_941));

	AOI22X1 i_82(
		.A0(n_793),
		.A1(n_787),
		.B0(n_7200),
		.B1(n_802),
		.Y(n_943));

	AOI221XL i_430(
		.A0(n_835),
		.A1(n_485),
		.B0(ir[9]),
		.B1(n_836),
		.C0(n_584),
		.Y(n_945));

	NOR2X1 i_114(
		.A(n_859),
		.B(reset),
		.Y(n_948));

	NOR2BX1 i_435(
		.AN(n_1105),
		.B(n_493),
		.Y(n_949));

	NOR2BX1 i_138(
		.AN(n_382),
		.B(n_932),
		.Y(n_950));

	NAND2X1 i_184(
		.A(n_950),
		.B(n_864),
		.Y(n_951));

	NOR3X1 i_2136(
		.A(n_824),
		.B(n_7200),
		.C(n_790),
		.Y(n_952));

	SDFFRHQX1 branch_stall_delay_reg(
		.SI(update_stall),
		.SE(scan_en),
		.D(n_3104),
		.CK(clk),
		.RN(n_7035),
		.Q(branch_stall_delay));

	OAI21XL i_3342(
		.A0(n_2515),
		.A1(n_1103),
		.B0(n_3107),
		.Y(n_3104));

	NAND2X1 i_3344(
		.A(n_2515),
		.B(branch_stall_delay),
		.Y(n_3107));

	NOR2X1 i_139(
		.A(n_496),
		.B(n_952),
		.Y(n_954));

	SDFFRHQX1 branch_stall_reg(
		.SI(branch_stall_delay),
		.SE(scan_en),
		.D(n_3110),
		.CK(clk),
		.RN(n_7035),
		.Q(branch_stall));

	OAI31X1 i_3349(
		.A0(n_383),
		.A1(n_407),
		.A2(n_4083),
		.B0(n_3113),
		.Y(n_3110));

	NAND3X1 i_3352(
		.A(n_407),
		.B(branch_stall),
		.C(n_1103),
		.Y(n_3113));

	NAND2BX1 i_442(
		.AN(n_704),
		.B(n_890),
		.Y(n_955));

	SDFFRHQX1 update_stall_reg(
		.SI(skip_one),
		.SE(scan_en),
		.D(n_3116),
		.CK(clk),
		.RN(n_7035),
		.Q(update_stall));

	MX2X1 i_3357(
		.S0(phi_1),
		.B(branch_stall),
		.A(update_stall),
		.Y(n_3116));

	SDFFRHQX1 three_cycle_reg(
		.SI(go_port),
		.SE(scan_en),
		.D(n_3122),
		.CK(clk),
		.RN(n_7035),
		.Q(SPCASCAN_N35_three_cycle));

	MX2X1 i_3364(
		.S0(n_2765),
		.B(n_2768),
		.A(SPCASCAN_N35_three_cycle),
		.Y(n_3122));

	SDFFRHQX1 two_cycle_reg(
		.SI(dmov_inc),
		.SE(scan_en),
		.D(n_4093),
		.CK(clk),
		.RN(n_7035),
		.Q(SPCASCAN_N32_two_cycle));

	AOI21X1 i_3371(
		.A0(n_1833),
		.A1(SPCASCAN_N32_two_cycle),
		.B0(n_3130),
		.Y(n_3128));

	AOI31X1 i_3372(
		.A0(n_1114),
		.A1(n_1062),
		.A2(n_1111),
		.B0(n_1833),
		.Y(n_3130));

	SDFFRHQX1 update_it_reg(
		.SI(branch_stall),
		.SE(scan_en),
		.D(n_3134),
		.CK(clk),
		.RN(n_4221),
		.Q(update_it));

	OAI21XL i_3378(
		.A0(n_1105),
		.A1(n_3146),
		.B0(n_3137),
		.Y(n_3134));

	NAND2X1 i_3380(
		.A(n_3146),
		.B(update_it),
		.Y(n_3137));

	NAND2X1 i_48(
		.A(phi_3),
		.B(n_4076),
		.Y(n_959));

	SDFFHQX1 acc_reg_0(
		.SI(acc[14]),
		.SE(scan_en),
		.D(n_3140),
		.CK(clk),
		.Q(acc[0]));

	OAI2BB1X1 i_3385(
		.A0N(n_4094),
		.A1N(acc[0]),
		.B0(n_3142),
		.Y(n_3140));

	NAND2X1 i_3386(
		.A(alu_result[0]),
		.B(\nbus_440[0] ),
		.Y(n_3142));

	NOR2X1 i_449(
		.A(n_959),
		.B(n_4077),
		.Y(n_960));

	SEDFFX1 acc_reg_1(
		.SI(acc[5]),
		.SE(scan_en),
		.D(alu_result[1]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[1]));

	SEDFFX1 acc_reg_2(
		.SI(top[15]),
		.SE(scan_en),
		.D(alu_result[2]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[2]));

	NOR2X1 i_135(
		.A(n_952),
		.B(n_584),
		.Y(n_962));

	SEDFFX1 acc_reg_3(
		.SI(pc[12]),
		.SE(scan_en),
		.D(alu_result[3]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[3]));

	SEDFFX1 acc_reg_4(
		.SI(acc[7]),
		.SE(scan_en),
		.D(alu_result[4]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[4]));

	SEDFFX1 acc_reg_5(
		.SI(acc[6]),
		.SE(scan_en),
		.D(alu_result[5]),
		.CK(clk),
		.E(\nbus_440[0] ),
		.Q(acc[5]));

	NAND2X1 i_140(
		.A(pc[11]),
		.B(pc[14]),
		.Y(n_965));

	SEDFFX1 acc_reg_6(
		.SI(acc[4]),
		.SE(scan_en),
		.D(alu_result[6]),
		.CK(clk),
		.E(\nbus_440[0] ),
		.Q(acc[6]));

	NAND2X1 i_1(
		.A(pc[0]),
		.B(pc[1]),
		.Y(n_966));

	SEDFFX1 acc_reg_7(
		.SI(acc[3]),
		.SE(scan_en),
		.D(alu_result[7]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[7]));

	NAND3X1 i_58(
		.A(pc[0]),
		.B(pc[1]),
		.C(pc[2]),
		.Y(n_967));

	SEDFFX1 acc_reg_8(
		.SI(acc[11]),
		.SE(scan_en),
		.D(alu_result[8]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[8]));

	NAND2BX1 i_108(
		.AN(n_967),
		.B(pc[3]),
		.Y(n_968));

	SEDFFX1 acc_reg_9(
		.SI(n_7862),
		.SE(scan_en),
		.D(alu_result[9]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[9]));

	NAND2BX1 i_361755(
		.AN(n_968),
		.B(pc[4]),
		.Y(n_969));

	SEDFFX1 acc_reg_10(
		.SI(acc[9]),
		.SE(scan_en),
		.D(alu_result[10]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[10]));

	NAND2BX1 i_56(
		.AN(n_969),
		.B(pc[5]),
		.Y(n_970));

	SEDFFX1 acc_reg_11(
		.SI(acc[10]),
		.SE(scan_en),
		.D(alu_result[11]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[11]));

	NAND2BX1 i_107(
		.AN(n_970),
		.B(pc[6]),
		.Y(n_971));

	SEDFFX1 acc_reg_12(
		.SI(acc[13]),
		.SE(scan_en),
		.D(alu_result[12]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[12]));

	NAND2BX1 i_30(
		.AN(n_971),
		.B(pc[7]),
		.Y(n_972));

	SEDFFX1 acc_reg_13(
		.SI(acc[8]),
		.SE(scan_en),
		.D(alu_result[13]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[13]));

	NAND2BX1 i_143(
		.AN(n_972),
		.B(pc[8]),
		.Y(n_973));

	SEDFFX1 acc_reg_14(
		.SI(read_prog),
		.SE(scan_en),
		.D(alu_result[14]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[14]));

	NAND2BX1 i_57(
		.AN(n_973),
		.B(pc[9]),
		.Y(n_974));

	SEDFFX1 acc_reg_15(
		.SI(acc[12]),
		.SE(scan_en),
		.D(alu_result[15]),
		.CK(clk),
		.E(n_7384),
		.Q(acc[15]));

	NAND2BX1 i_581765(
		.AN(n_974),
		.B(pc[10]),
		.Y(n_975));

	SEDFFX1 acc_reg_16(
		.SI(acc[18]),
		.SE(scan_en),
		.D(alu_result[16]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[16]));

	NAND2X1 i_68(
		.A(pc[13]),
		.B(pc[12]),
		.Y(n_976));

	SEDFFX1 acc_reg_17(
		.SI(acc[0]),
		.SE(scan_en),
		.D(alu_result[17]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[17]));

	SEDFFX1 acc_reg_18(
		.SI(acc[17]),
		.SE(scan_en),
		.D(alu_result[18]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[18]));

	NOR3X1 i_159(
		.A(n_975),
		.B(n_976),
		.C(n_965),
		.Y(n_978));

	SEDFFX1 acc_reg_19(
		.SI(acc[22]),
		.SE(scan_en),
		.D(alu_result[19]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[19]));

	NAND2X1 i_42(
		.A(pc[10]),
		.B(pc[11]),
		.Y(n_979));

	SEDFFX1 acc_reg_20(
		.SI(acc[23]),
		.SE(scan_en),
		.D(alu_result[20]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[20]));

	SEDFFX1 acc_reg_21(
		.SI(acc[24]),
		.SE(scan_en),
		.D(alu_result[21]),
		.CK(clk),
		.E(\nbus_440[0] ),
		.Q(acc[21]));

	NOR3X1 i_156(
		.A(n_979),
		.B(n_976),
		.C(n_974),
		.Y(n_981));

	SEDFFX1 acc_reg_22(
		.SI(SPCASCAN_N36_tdsp_state_1_),
		.SE(scan_en),
		.D(alu_result[22]),
		.CK(clk),
		.E(\nbus_440[0] ),
		.Q(acc[22]));

	NAND3X1 i_69(
		.A(pc[10]),
		.B(pc[11]),
		.C(pc[9]),
		.Y(n_982));

	SEDFFX1 acc_reg_23(
		.SI(acc[16]),
		.SE(scan_en),
		.D(alu_result[23]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[23]));

	SEDFFX1 acc_reg_24(
		.SI(SPCASCAN_N33_samp_int),
		.SE(scan_en),
		.D(alu_result[24]),
		.CK(clk),
		.E(\nbus_440[0] ),
		.Q(acc[24]));

	NOR3X1 i_157(
		.A(n_973),
		.B(n_982),
		.C(n_4101),
		.Y(n_984));

	SEDFFX1 acc_reg_25(
		.SI(acc[30]),
		.SE(scan_en),
		.D(alu_result[25]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[25]));

	SEDFFX1 acc_reg_26(
		.SI(acc[25]),
		.SE(scan_en),
		.D(alu_result[26]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[26]));

	SEDFFX1 acc_reg_27(
		.SI(acc[28]),
		.SE(scan_en),
		.D(alu_result[27]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[27]));

	SEDFFX1 acc_reg_28(
		.SI(acc[26]),
		.SE(scan_en),
		.D(alu_result[28]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[28]));

	SEDFFX1 acc_reg_29(
		.SI(acc[31]),
		.SE(scan_en),
		.D(alu_result[29]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[29]));

	NAND3X1 i_155(
		.A(n_926),
		.B(n_886),
		.C(n_4080),
		.Y(n_989));

	SEDFFX1 acc_reg_30(
		.SI(SPCASCAN_N31_tdsp_state_2_),
		.SE(scan_en),
		.D(alu_result[30]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[30]));

	SEDFFX1 acc_reg_31(
		.SI(acc[27]),
		.SE(scan_en),
		.D(alu_result[31]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[31]));

	SEDFFX1 acc_reg_32(
		.SI(acc[29]),
		.SE(scan_en),
		.D(alu_result[32]),
		.CK(clk),
		.E(n_7353),
		.Q(acc[32]));

	NAND3BX1 i_13(
		.AN(arp),
		.B(n_876),
		.C(n_1105),
		.Y(n_992));

	SDFFRHQX1 arp_reg(
		.SI(sel_op_b[1]),
		.SE(scan_en),
		.D(n_3340),
		.CK(clk),
		.RN(n_4221),
		.Q(arp));

	OAI2BB1X1 i_3621(
		.A0N(ir[0]),
		.A1N(n_1104),
		.B0(n_3343),
		.Y(n_3340));

	NAND2BX1 i_3623(
		.AN(n_1104),
		.B(arp),
		.Y(n_3343));

	SDFFHQX1 null_op_reg0(
		.SI(ar1[3]),
		.SE(scan_en),
		.D(n_3349),
		.CK(clk),
		.Q(Q));

	AND2X1 i_3630(
		.A(n_2909),
		.B(Q),
		.Y(n_3349));

	OR3XL i_65(
		.A(ar[0]),
		.B(ar[1]),
		.C(ar[2]),
		.Y(n_994));

	SDFFRHQX1 ovm_reg(
		.SI(update_it),
		.SE(scan_en),
		.D(n_3352),
		.CK(clk),
		.RN(n_4221),
		.Q(ovm));

	OAI21XL i_3635(
		.A0(n_1108),
		.A1(n_4223),
		.B0(n_3354),
		.Y(n_3352));

	NAND4BXL i_3636(
		.AN(ir[2]),
		.B(ir[0]),
		.C(n_1108),
		.D(n_869),
		.Y(n_3354));

	NOR2X1 i_98(
		.A(n_994),
		.B(ar[3]),
		.Y(n_995));

	SEDFFX1 sel_op_b_reg_0(
		.SI(sel_op_a[2]),
		.SE(scan_en),
		.D(nbus_439[0]),
		.CK(clk),
		.E(\nbus_434[0] ),
		.Q(sel_op_b[0]));

	NOR2X1 i_129(
		.A(n_4074),
		.B(ar[4]),
		.Y(n_996));

	SEDFFX1 sel_op_b_reg_1(
		.SI(sel_op_b[2]),
		.SE(scan_en),
		.D(nbus_439[1]),
		.CK(clk),
		.E(\nbus_434[0] ),
		.Q(sel_op_b[1]));

	OR3XL i_130(
		.A(ar[4]),
		.B(ar[5]),
		.C(n_4074),
		.Y(n_997));

	SEDFFX1 sel_op_b_reg_2(
		.SI(sel_op_a[0]),
		.SE(scan_en),
		.D(nbus_439[2]),
		.CK(clk),
		.E(\nbus_434[0] ),
		.Q(sel_op_b[2]));

	NOR2X1 i_131(
		.A(n_997),
		.B(ar[6]),
		.Y(n_998));

	SDFFRHQX1 skip_one_reg(
		.SI(acc[32]),
		.SE(scan_en),
		.D(n_3376),
		.CK(clk),
		.RN(n_4221),
		.Q(skip_one));

	OAI21XL i_3664(
		.A0(n_1793),
		.A1(n_1790),
		.B0(n_3379),
		.Y(n_3376));

	NAND2X1 i_3666(
		.A(n_1790),
		.B(skip_one),
		.Y(n_3379));

	NOR2X1 i_34(
		.A(n_4073),
		.B(ar[7]),
		.Y(n_999));

	SDFFRHQX1 ov_flag_reg(
		.SI(ovm),
		.SE(scan_en),
		.D(n_3382),
		.CK(clk),
		.RN(n_4221),
		.Q(SPCASCAN_N30_ov));

	OAI21XL i_3671(
		.A0(n_2387),
		.A1(n_2384),
		.B0(n_3385),
		.Y(n_3382));

	NAND2X1 i_3673(
		.A(n_2384),
		.B(SPCASCAN_N30_ov),
		.Y(n_3385));

	OR3XL i_163(
		.A(ar[7]),
		.B(ar[8]),
		.C(n_4073),
		.Y(n_1000));

	SDFFSHQX1 pc_reg_0(
		.SI(pc[2]),
		.SE(scan_en),
		.D(n_3388),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[0]));

	MX2X1 i_3678(
		.S0(n_7513),
		.B(nbus_437[0]),
		.A(pc[0]),
		.Y(n_3388));

	NOR2X1 i_164(
		.A(n_1000),
		.B(ar[9]),
		.Y(n_1001));

	SDFFSHQX1 pc_reg_1(
		.SI(FE_PT1_),
		.SE(scan_en),
		.D(n_3394),
		.CK(clk),
		.SN(n_4221),
		.Q(pc[1]));

	MX2X1 i_3685(
		.S0(n_7513),
		.B(nbus_437[1]),
		.A(pc[1]),
		.Y(n_3394));

	NOR2X1 i_165(
		.A(n_4072),
		.B(ar[10]),
		.Y(n_1002));

	SDFFSHQX1 pc_reg_2(
		.SI(SPCASCAN_N23_done),
		.SE(scan_en),
		.D(n_3400),
		.CK(clk),
		.SN(n_4221),
		.Q(pc[2]));

	MX2X1 i_3692(
		.S0(n_7513),
		.B(nbus_437[2]),
		.A(pc[2]),
		.Y(n_3400));

	SDFFSHQX1 pc_reg_3(
		.SI(decode[4]),
		.SE(scan_en),
		.D(n_3406),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[3]));

	MX2X1 i_3699(
		.S0(n_7513),
		.B(nbus_437[3]),
		.A(pc[3]),
		.Y(n_3406));

	SDFFSHQX1 pc_reg_4(
		.SI(decode[6]),
		.SE(scan_en),
		.D(n_3412),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[4]));

	MX2X1 i_3706(
		.S0(n_7513),
		.B(nbus_437[4]),
		.A(pc[4]),
		.Y(n_3412));

	NOR4X1 i_566(
		.A(ar[11]),
		.B(ar[12]),
		.C(ar[13]),
		.D(ar[14]),
		.Y(n_1005));

	SDFFSHQX1 pc_reg_5(
		.SI(p[17]),
		.SE(scan_en),
		.D(n_3418),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[5]));

	MX2X1 i_3713(
		.S0(n_7513),
		.B(nbus_437[5]),
		.A(pc[5]),
		.Y(n_3418));

	NAND2X1 i_169(
		.A(n_1002),
		.B(n_1005),
		.Y(n_1006));

	SDFFSHQX1 pc_reg_6(
		.SI(pc[5]),
		.SE(scan_en),
		.D(n_3424),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[6]));

	MX2X1 i_3720(
		.S0(n_7513),
		.B(nbus_437[6]),
		.A(pc[6]),
		.Y(n_3424));

	SDFFSHQX1 pc_reg_7(
		.SI(pc[6]),
		.SE(scan_en),
		.D(n_3430),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[7]));

	MX2X1 i_3727(
		.S0(n_7513),
		.B(nbus_437[7]),
		.A(pc[7]),
		.Y(n_3430));

	NAND3BX1 i_12(
		.AN(arp),
		.B(n_908),
		.C(n_1105),
		.Y(n_1008));

	SDFFSHQX1 pc_reg_8(
		.SI(decode[2]),
		.SE(scan_en),
		.D(n_3436),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[8]));

	MX2X1 i_3735(
		.S0(n_7513),
		.B(nbus_437[8]),
		.A(pc[8]),
		.Y(n_3436));

	NAND2X1 i_12042(
		.A(ar[0]),
		.B(ar[1]),
		.Y(n_1009));

	SDFFSHQX1 pc_reg_9(
		.SI(acc[2]),
		.SE(scan_en),
		.D(n_3442),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[9]));

	MX2X1 i_3743(
		.S0(n_7513),
		.B(nbus_437[9]),
		.A(pc[9]),
		.Y(n_3442));

	NAND3X1 i_64(
		.A(ar[0]),
		.B(ar[1]),
		.C(ar[2]),
		.Y(n_1010));

	SDFFSHQX1 pc_reg_10(
		.SI(pc[11]),
		.SE(scan_en),
		.D(n_3448),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[10]));

	MX2X1 i_3751(
		.S0(\nbus_436[0] ),
		.B(nbus_437[10]),
		.A(pc[10]),
		.Y(n_3448));

	NAND2BX1 i_192059(
		.AN(n_1010),
		.B(ar[3]),
		.Y(n_1011));

	SDFFSHQX1 pc_reg_11(
		.SI(pc[15]),
		.SE(scan_en),
		.D(n_3454),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[11]));

	MX2X1 i_3758(
		.S0(n_7513),
		.B(nbus_437[11]),
		.A(pc[11]),
		.Y(n_3454));

	NAND2BX1 i_59(
		.AN(n_1011),
		.B(ar[4]),
		.Y(n_1012));

	SDFFSHQX1 pc_reg_12(
		.SI(pc[9]),
		.SE(scan_en),
		.D(n_3460),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[12]));

	MXI2X1 i_3765(
		.S0(n_7513),
		.B(nbus_437[12]),
		.A(n_4101),
		.Y(n_3460));

	NAND2BX1 i_372075(
		.AN(n_1012),
		.B(ar[5]),
		.Y(n_1013));

	SDFFSHQX1 pc_reg_13(
		.SI(dec_go_data),
		.SE(scan_en),
		.D(n_3466),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[13]));

	MX2X1 i_3772(
		.S0(n_7513),
		.B(nbus_437[13]),
		.A(pc[13]),
		.Y(n_3466));

	NAND2BX1 i_382076(
		.AN(n_1013),
		.B(ar[6]),
		.Y(n_1014));

	SDFFSHQX1 pc_reg_14(
		.SI(pc[13]),
		.SE(scan_en),
		.D(n_3472),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[14]));

	MX2X1 i_3779(
		.S0(n_7513),
		.B(nbus_437[14]),
		.A(pc[14]),
		.Y(n_3472));

	NAND2BX1 i_53(
		.AN(n_1014),
		.B(ar[7]),
		.Y(n_1015));

	SDFFSHQX1 pc_reg_15(
		.SI(pc[14]),
		.SE(scan_en),
		.D(n_3478),
		.CK(clk),
		.SN(n_6303),
		.Q(pc[15]));

	MX2X1 i_3786(
		.S0(n_7513),
		.B(nbus_437[15]),
		.A(pc[15]),
		.Y(n_3478));

	SDFFRHQX1 read_prog_reg(
		.SI(go_prog),
		.SE(scan_en),
		.D(n_3484),
		.CK(clk),
		.RN(n_7035),
		.Q(read_prog));

	OAI21XL i_3793(
		.A0(n_2610),
		.A1(n_1940),
		.B0(n_3487),
		.Y(n_3484));

	NAND2X1 i_3795(
		.A(n_1940),
		.B(read_prog),
		.Y(n_3487));

	NAND3BX1 i_191(
		.AN(n_1015),
		.B(ar[9]),
		.C(ar[8]),
		.Y(n_1017));

	SDFFRHQX1 dp_reg(
		.SI(sel_op_a[1]),
		.SE(scan_en),
		.D(n_3490),
		.CK(clk),
		.RN(n_7035),
		.Q(dp));

	OAI21XL i_3800(
		.A0(n_2534),
		.A1(n_1107),
		.B0(n_3493),
		.Y(n_3490));

	NAND2X1 i_3802(
		.A(n_1107),
		.B(dp),
		.Y(n_3493));

	NAND2BX1 i_582093(
		.AN(n_1017),
		.B(ar[10]),
		.Y(n_1018));

	SEDFFX1 sel_op_a_reg_0(
		.SI(dec_go_port),
		.SE(scan_en),
		.D(nbus_435[0]),
		.CK(clk),
		.E(\nbus_434[0] ),
		.Q(sel_op_a[0]));

	SEDFFX1 sel_op_a_reg_1(
		.SI(sel_op_b[0]),
		.SE(scan_en),
		.D(nbus_435[1]),
		.CK(clk),
		.E(\nbus_434[0] ),
		.Q(sel_op_a[1]));

	SEDFFX1 sel_op_a_reg_2(
		.SI(Q),
		.SE(scan_en),
		.D(nbus_435[2]),
		.CK(clk),
		.E(\nbus_434[0] ),
		.Q(sel_op_a[2]));

	NAND4X1 i_561(
		.A(ar[11]),
		.B(ar[12]),
		.C(ar[14]),
		.D(ar[13]),
		.Y(n_1021));

	SDFFRHQX1 go_port_reg(
		.SI(phi_5),
		.SE(scan_en),
		.D(n_3514),
		.CK(clk),
		.RN(n_7035),
		.Q(go_port));

	OAI31X1 i_3828(
		.A0(n_830),
		.A1(n_2115),
		.A2(n_832),
		.B0(n_3517),
		.Y(n_3514));

	NAND2X1 i_3830(
		.A(n_2115),
		.B(go_port),
		.Y(n_3517));

	NOR2X1 i_622097(
		.A(n_1018),
		.B(n_1021),
		.Y(n_1022));

	SEDFFX1 top_reg_0(
		.SI(top[14]),
		.SE(scan_en),
		.D(mdr[0]),
		.CK(clk),
		.E(n_6809),
		.Q(top[0]));

	SEDFFX1 top_reg_1(
		.SI(top[6]),
		.SE(scan_en),
		.D(mdr[1]),
		.CK(clk),
		.E(n_6809),
		.Q(top[1]));

	SEDFFX1 top_reg_2(
		.SI(top[7]),
		.SE(scan_en),
		.D(mdr[2]),
		.CK(clk),
		.E(n_6809),
		.Q(top[2]));

	OR3XL i_166(
		.A(ar[10]),
		.B(ar[11]),
		.C(n_4072),
		.Y(n_1025));

	SEDFFX1 top_reg_3(
		.SI(top[2]),
		.SE(scan_en),
		.D(mdr[3]),
		.CK(clk),
		.E(n_6809),
		.Q(top[3]));

	NOR2X1 i_167(
		.A(ar[12]),
		.B(n_1025),
		.Y(n_1026));

	SEDFFX1 top_reg_4(
		.SI(top[5]),
		.SE(scan_en),
		.D(mdr[4]),
		.CK(clk),
		.E(\nbus_432[0] ),
		.Q(top[4]));

	NOR2X1 i_168(
		.A(n_4075),
		.B(ar[13]),
		.Y(n_1027));

	SEDFFX1 top_reg_5(
		.SI(top[12]),
		.SE(scan_en),
		.D(mdr[5]),
		.CK(clk),
		.E(\nbus_432[0] ),
		.Q(top[5]));

	NAND2X1 i_197(
		.A(ar[11]),
		.B(ar[10]),
		.Y(n_1028));

	SEDFFX1 top_reg_6(
		.SI(top[9]),
		.SE(scan_en),
		.D(mdr[6]),
		.CK(clk),
		.E(n_6809),
		.Q(top[6]));

	NOR2X1 i_592094(
		.A(n_1017),
		.B(n_1028),
		.Y(n_1029));

	SEDFFX1 top_reg_7(
		.SI(top[4]),
		.SE(scan_en),
		.D(mdr[7]),
		.CK(clk),
		.E(\nbus_432[0] ),
		.Q(top[7]));

	SEDFFX1 top_reg_8(
		.SI(ir[1]),
		.SE(scan_en),
		.D(mdr[8]),
		.CK(clk),
		.E(n_6809),
		.Q(top[8]));

	NAND3X1 i_612096(
		.A(ar[13]),
		.B(ar[12]),
		.C(n_1029),
		.Y(n_1031));

	SEDFFX1 top_reg_9(
		.SI(top[13]),
		.SE(scan_en),
		.D(mdr[9]),
		.CK(clk),
		.E(n_6809),
		.Q(top[9]));

	SEDFFX1 top_reg_10(
		.SI(top[8]),
		.SE(scan_en),
		.D(mdr[10]),
		.CK(clk),
		.E(n_6809),
		.Q(top[10]));

	NAND2BX1 i_562091(
		.AN(n_1015),
		.B(ar[8]),
		.Y(n_1033));

	SEDFFX1 top_reg_11(
		.SI(top[10]),
		.SE(scan_en),
		.D(mdr[11]),
		.CK(clk),
		.E(n_6809),
		.Q(top[11]));

	SEDFFX1 top_reg_12(
		.SI(top[1]),
		.SE(scan_en),
		.D(mdr[12]),
		.CK(clk),
		.E(n_6809),
		.Q(top[12]));

	NAND4X1 i_585(
		.A(ar[11]),
		.B(ar[10]),
		.C(ar[12]),
		.D(ar[9]),
		.Y(n_1035));

	SEDFFX1 top_reg_13(
		.SI(top[0]),
		.SE(scan_en),
		.D(mdr[13]),
		.CK(clk),
		.E(n_6809),
		.Q(top[13]));

	OR2X1 i_602095(
		.A(n_1033),
		.B(n_1035),
		.Y(n_1036));

	SEDFFX1 top_reg_14(
		.SI(acc[1]),
		.SE(scan_en),
		.D(mdr[14]),
		.CK(clk),
		.E(n_6809),
		.Q(top[14]));

	SEDFFX1 top_reg_15(
		.SI(ir[12]),
		.SE(scan_en),
		.D(mdr[15]),
		.CK(clk),
		.E(n_6809),
		.Q(top[15]));

	SDFFRHQX1 dmov_inc_reg(
		.SI(phi_1),
		.SE(scan_en),
		.D(n_3616),
		.CK(clk),
		.RN(n_7035),
		.Q(dmov_inc));

	MX2X1 i_3949(
		.S0(n_2235),
		.B(n_4081),
		.A(dmov_inc),
		.Y(n_3616));

	SDFFRHQX1 read_data_reg(
		.SI(phi_3),
		.SE(scan_en),
		.D(n_3625),
		.CK(clk),
		.RN(n_7035),
		.Q(read_data));

	AND2X1 i_3958(
		.A(n_2079),
		.B(read_data),
		.Y(n_3625));

	SDFFRHQX1 read_port_reg(
		.SI(n_7866),
		.SE(scan_en),
		.D(n_3631),
		.CK(clk),
		.RN(n_7035),
		.Q(read_port));

	AND2X1 i_3966(
		.A(n_2115),
		.B(read_port),
		.Y(n_3631));

	SDFFRHQX1 go_data_reg(
		.SI(dec_go_prog),
		.SE(scan_en),
		.D(n_3634),
		.CK(clk),
		.RN(n_7035),
		.Q(go_data));

	OAI21XL i_3971(
		.A0(n_2079),
		.A1(n_2082),
		.B0(n_3637),
		.Y(n_3634));

	NAND2X1 i_3973(
		.A(n_2079),
		.B(go_data),
		.Y(n_3637));

	SEDFFX1 ar0_reg_0(
		.SI(ar1[1]),
		.SE(scan_en),
		.D(nbus_431[0]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[0]));

	NOR2X1 i_16(
		.A(n_1105),
		.B(n_824),
		.Y(n_1043));

	SEDFFX1 ar0_reg_1(
		.SI(ar1[13]),
		.SE(scan_en),
		.D(nbus_431[1]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[1]));

	AOI22X1 i_144(
		.A0(ir[7]),
		.A1(n_1043),
		.B0(mdr[7]),
		.B1(n_7029),
		.Y(n_1044));

	SEDFFX1 ar0_reg_2(
		.SI(port_as),
		.SE(scan_en),
		.D(nbus_431[2]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[2]));

	AOI2BB1X1 i_642(
		.A0N(n_751),
		.A1N(n_7203),
		.B0(n_644),
		.Y(n_1045));

	SEDFFX1 ar0_reg_3(
		.SI(ar1[2]),
		.SE(scan_en),
		.D(nbus_431[3]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[3]));

	AOI22X1 i_145(
		.A0(ir[6]),
		.A1(n_1043),
		.B0(mdr[6]),
		.B1(n_7029),
		.Y(n_1046));

	SEDFFX1 ar0_reg_4(
		.SI(ar1[4]),
		.SE(scan_en),
		.D(nbus_431[4]),
		.CK(clk),
		.E(\nbus_430[0] ),
		.Q(ar0[4]));

	AOI2BB1X1 i_651(
		.A0N(n_755),
		.A1N(n_7203),
		.B0(n_651),
		.Y(n_1047));

	SEDFFX1 ar0_reg_5(
		.SI(ar1[7]),
		.SE(scan_en),
		.D(nbus_431[5]),
		.CK(clk),
		.E(\nbus_430[0] ),
		.Q(ar0[5]));

	AOI22X1 i_146(
		.A0(ir[5]),
		.A1(n_1043),
		.B0(mdr[5]),
		.B1(n_7029),
		.Y(n_1048));

	SEDFFX1 ar0_reg_6(
		.SI(ar1[6]),
		.SE(scan_en),
		.D(nbus_431[6]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[6]));

	AOI2BB1X1 i_660(
		.A0N(n_759),
		.A1N(n_7206),
		.B0(n_658),
		.Y(n_1049));

	SEDFFX1 ar0_reg_7(
		.SI(ar1[5]),
		.SE(scan_en),
		.D(nbus_431[7]),
		.CK(clk),
		.E(\nbus_430[0] ),
		.Q(ar0[7]));

	AOI22X1 i_147(
		.A0(ir[4]),
		.A1(n_1043),
		.B0(mdr[4]),
		.B1(n_7029),
		.Y(n_1050));

	SEDFFX1 ar0_reg_8(
		.SI(ar1[8]),
		.SE(scan_en),
		.D(nbus_431[8]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[8]));

	AOI2BB1X1 i_669(
		.A0N(n_763),
		.A1N(n_7203),
		.B0(n_665),
		.Y(n_1051));

	SEDFFX1 ar0_reg_9(
		.SI(ar0[12]),
		.SE(scan_en),
		.D(nbus_431[9]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[9]));

	AOI22X1 i_148(
		.A0(ir[3]),
		.A1(n_1043),
		.B0(mdr[3]),
		.B1(n_7029),
		.Y(n_1052));

	SEDFFX1 ar0_reg_10(
		.SI(ar0[9]),
		.SE(scan_en),
		.D(nbus_431[10]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[10]));

	AOI2BB1X1 i_678(
		.A0N(n_767),
		.A1N(n_7203),
		.B0(n_672),
		.Y(n_1053));

	SEDFFX1 ar0_reg_11(
		.SI(ar1[10]),
		.SE(scan_en),
		.D(nbus_431[11]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[11]));

	AOI22X1 i_149(
		.A0(ir[2]),
		.A1(n_1043),
		.B0(mdr[2]),
		.B1(n_7029),
		.Y(n_1054));

	SEDFFX1 ar0_reg_12(
		.SI(ar1[12]),
		.SE(scan_en),
		.D(nbus_431[12]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[12]));

	AOI2BB1X1 i_687(
		.A0N(n_771),
		.A1N(n_7203),
		.B0(n_679),
		.Y(n_1055));

	SEDFFX1 ar0_reg_13(
		.SI(ar0[1]),
		.SE(scan_en),
		.D(nbus_431[13]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[13]));

	AOI22X1 i_150(
		.A0(ir[1]),
		.A1(n_1043),
		.B0(mdr[1]),
		.B1(n_7029),
		.Y(n_1056));

	SEDFFX1 ar0_reg_14(
		.SI(FE_PT2_),
		.SE(scan_en),
		.D(nbus_431[14]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[14]));

	OAI21XL i_105(
		.A0(ar[0]),
		.A1(ar[1]),
		.B0(n_1009),
		.Y(n_1057));

	SEDFFX1 ar0_reg_15(
		.SI(decode[8]),
		.SE(scan_en),
		.D(nbus_431[15]),
		.CK(clk),
		.E(n_7021),
		.Q(ar0[15]));

	MX2X1 i_693(
		.S0(n_1057),
		.B(n_7203),
		.A(n_7206),
		.Y(n_1058));

	SDFFRHQX1 go_prog_reg(
		.SI(acc[15]),
		.SE(scan_en),
		.D(n_3736),
		.CK(clk),
		.RN(n_7035),
		.Q(go_prog));

	OAI21XL i_4092(
		.A0(n_1940),
		.A1(n_1943),
		.B0(n_3739),
		.Y(n_3736));

	NAND2X1 i_4094(
		.A(n_1940),
		.B(go_prog),
		.Y(n_3739));

	SDFFRHQX1 fetch_branch_reg(
		.SI(alu_cmd[3]),
		.SE(scan_en),
		.D(n_4095),
		.CK(clk),
		.RN(n_7035),
		.Q(fetch_branch));

	AOI31X1 i_4099(
		.A0(n_1103),
		.A1(n_407),
		.A2(fetch_branch),
		.B0(n_3744),
		.Y(n_3742));

	AOI211X1 i_4100(
		.A0(phi_1),
		.A1(branch_stall),
		.B0(n_444),
		.C0(n_407),
		.Y(n_3744));

	SDFFHQX1 alu_cmd_reg_0(
		.SI(fetch_branch),
		.SE(scan_en),
		.D(n_4096),
		.CK(clk),
		.Q(\nbus_682[0] ));

	AOI21X1 i_4106(
		.A0(\nbus_428[0] ),
		.A1(\nbus_682[0] ),
		.B0(n_3750),
		.Y(n_3748));

	AOI31X1 i_4107(
		.A0(n_934),
		.A1(n_879),
		.A2(n_1071),
		.B0(\nbus_428[0] ),
		.Y(n_3750));

	AOI22X1 i_151(
		.A0(ir[0]),
		.A1(n_1043),
		.B0(mdr[0]),
		.B1(n_7029),
		.Y(n_1061));

	SDFFHQX1 alu_cmd_reg_1(
		.SI(\nbus_682[0] ),
		.SE(scan_en),
		.D(n_3754),
		.CK(clk),
		.Q(\nbus_681[1] ));

	OAI21XL i_4113(
		.A0(\nbus_428[0] ),
		.A1(\nbus_429[1] ),
		.B0(n_3757),
		.Y(n_3754));

	NAND2X1 i_4115(
		.A(\nbus_428[0] ),
		.B(\nbus_681[1] ),
		.Y(n_3757));

	AOI22X1 i_710(
		.A0(n_784),
		.A1(n_4088),
		.B0(n_829),
		.B1(n_802),
		.Y(n_1062));

	SEDFFX1 alu_cmd_reg_2(
		.SI(\nbus_681[1] ),
		.SE(scan_en),
		.D(\nbus_429[2] ),
		.CK(clk),
		.E(n_4097),
		.Q(alu_cmd[2]));

	SDFFHQX1 alu_cmd_reg_3(
		.SI(FE_PT4_),
		.SE(scan_en),
		.D(n_3769),
		.CK(clk),
		.Q(alu_cmd[3]));

	AND2X1 i_4129(
		.A(alu_cmd[3]),
		.B(\nbus_428[0] ),
		.Y(n_3769));

	NAND2X1 i_714(
		.A(n_7218),
		.B(n_817),
		.Y(n_1064));

	SEDFFX1 p_reg_0(
		.SI(p[1]),
		.SE(scan_en),
		.D(mpy_result[0]),
		.CK(clk),
		.E(n_7423),
		.Q(p[0]));

	OAI21XL i_123(
		.A0(ir[14]),
		.A1(n_820),
		.B0(n_926),
		.Y(n_1065));

	SEDFFX1 p_reg_1(
		.SI(p[4]),
		.SE(scan_en),
		.D(mpy_result[1]),
		.CK(clk),
		.E(n_7423),
		.Q(p[1]));

	SEDFFX1 p_reg_2(
		.SI(p[8]),
		.SE(scan_en),
		.D(mpy_result[2]),
		.CK(clk),
		.E(n_7423),
		.Q(p[2]));

	SEDFFX1 p_reg_3(
		.SI(p[16]),
		.SE(scan_en),
		.D(mpy_result[3]),
		.CK(clk),
		.E(n_7423),
		.Q(p[3]));

	AOI211X1 i_730(
		.A0(n_7200),
		.A1(n_823),
		.B0(n_470),
		.C0(n_1065),
		.Y(n_1068));

	SEDFFX1 p_reg_4(
		.SI(p[3]),
		.SE(scan_en),
		.D(mpy_result[4]),
		.CK(clk),
		.E(\nbus_426[0] ),
		.Q(p[4]));

	SEDFFX1 p_reg_5(
		.SI(p[27]),
		.SE(scan_en),
		.D(mpy_result[5]),
		.CK(clk),
		.E(\nbus_426[0] ),
		.Q(p[5]));

	SEDFFX1 p_reg_6(
		.SI(p[12]),
		.SE(scan_en),
		.D(mpy_result[6]),
		.CK(clk),
		.E(n_7423),
		.Q(p[6]));

	NOR4BX1 i_733(
		.AN(n_1068),
		.B(n_704),
		.C(n_467),
		.D(n_705),
		.Y(n_1071));

	SEDFFX1 p_reg_7(
		.SI(p[13]),
		.SE(scan_en),
		.D(mpy_result[7]),
		.CK(clk),
		.E(n_7423),
		.Q(p[7]));

	SEDFFX1 p_reg_8(
		.SI(p[14]),
		.SE(scan_en),
		.D(mpy_result[8]),
		.CK(clk),
		.E(n_7423),
		.Q(p[8]));

	SEDFFX1 p_reg_9(
		.SI(p[2]),
		.SE(scan_en),
		.D(mpy_result[9]),
		.CK(clk),
		.E(n_7423),
		.Q(p[9]));

	SEDFFX1 p_reg_10(
		.SI(p[15]),
		.SE(scan_en),
		.D(mpy_result[10]),
		.CK(clk),
		.E(n_7423),
		.Q(p[10]));

	SEDFFX1 p_reg_11(
		.SI(p[9]),
		.SE(scan_en),
		.D(mpy_result[11]),
		.CK(clk),
		.E(n_7423),
		.Q(p[11]));

	NAND4BXL i_753(
		.AN(n_812),
		.B(n_871),
		.C(n_790),
		.D(n_713),
		.Y(n_1076));

	SEDFFX1 p_reg_12(
		.SI(p[7]),
		.SE(scan_en),
		.D(mpy_result[12]),
		.CK(clk),
		.E(n_7423),
		.Q(p[12]));

	SEDFFX1 p_reg_13(
		.SI(p[0]),
		.SE(scan_en),
		.D(mpy_result[13]),
		.CK(clk),
		.E(n_7423),
		.Q(p[13]));

	SEDFFX1 p_reg_14(
		.SI(p[10]),
		.SE(scan_en),
		.D(mpy_result[14]),
		.CK(clk),
		.E(n_7423),
		.Q(p[14]));

	SEDFFX1 p_reg_15(
		.SI(p[6]),
		.SE(scan_en),
		.D(mpy_result[15]),
		.CK(clk),
		.E(n_7423),
		.Q(p[15]));

	SEDFFX1 p_reg_16(
		.SI(p[21]),
		.SE(scan_en),
		.D(mpy_result[16]),
		.CK(clk),
		.E(n_6812),
		.Q(p[16]));

	NAND4X1 i_756(
		.A(n_715),
		.B(n_714),
		.C(n_943),
		.D(n_716),
		.Y(n_1081));

	SEDFFX1 p_reg_17(
		.SI(p[11]),
		.SE(scan_en),
		.D(mpy_result[17]),
		.CK(clk),
		.E(n_6812),
		.Q(p[17]));

	SEDFFX1 p_reg_18(
		.SI(p[28]),
		.SE(scan_en),
		.D(mpy_result[18]),
		.CK(clk),
		.E(n_6812),
		.Q(p[18]));

	SEDFFX1 p_reg_19(
		.SI(p[20]),
		.SE(scan_en),
		.D(mpy_result[19]),
		.CK(clk),
		.E(n_6812),
		.Q(p[19]));

	NAND3X1 i_159005(
		.A(arp),
		.B(n_876),
		.C(n_1105),
		.Y(n_1084));

	SEDFFX1 p_reg_20(
		.SI(p[22]),
		.SE(scan_en),
		.D(mpy_result[20]),
		.CK(clk),
		.E(n_6812),
		.Q(p[20]));

	SEDFFX1 p_reg_21(
		.SI(p[30]),
		.SE(scan_en),
		.D(mpy_result[21]),
		.CK(clk),
		.E(n_6812),
		.Q(p[21]));

	NAND3X1 i_14(
		.A(arp),
		.B(n_1105),
		.C(n_908),
		.Y(n_1086));

	SEDFFX1 p_reg_22(
		.SI(SPCASCAN_N7_present_state_1_),
		.SE(scan_en),
		.D(mpy_result[22]),
		.CK(clk),
		.E(n_6812),
		.Q(p[22]));

	SEDFFX1 p_reg_23(
		.SI(p[19]),
		.SE(scan_en),
		.D(mpy_result[23]),
		.CK(clk),
		.E(n_6812),
		.Q(p[23]));

	SEDFFX1 p_reg_24(
		.SI(p[18]),
		.SE(scan_en),
		.D(mpy_result[24]),
		.CK(clk),
		.E(n_6812),
		.Q(p[24]));

	SEDFFX1 p_reg_25(
		.SI(p[23]),
		.SE(scan_en),
		.D(mpy_result[25]),
		.CK(clk),
		.E(n_6812),
		.Q(p[25]));

	SEDFFX1 p_reg_26(
		.SI(ir[6]),
		.SE(scan_en),
		.D(mpy_result[26]),
		.CK(clk),
		.E(\nbus_426[0] ),
		.Q(p[26]));

	SEDFFX1 p_reg_27(
		.SI(p[26]),
		.SE(scan_en),
		.D(mpy_result[27]),
		.CK(clk),
		.E(\nbus_426[0] ),
		.Q(p[27]));

	SEDFFX1 p_reg_28(
		.SI(SPCASCAN_N6_present_state_2_),
		.SE(scan_en),
		.D(mpy_result[28]),
		.CK(clk),
		.E(n_6812),
		.Q(p[28]));

	SEDFFX1 p_reg_29(
		.SI(p[31]),
		.SE(scan_en),
		.D(mpy_result[29]),
		.CK(clk),
		.E(n_6812),
		.Q(p[29]));

	SEDFFX1 p_reg_30(
		.SI(p[5]),
		.SE(scan_en),
		.D(mpy_result[30]),
		.CK(clk),
		.E(n_6812),
		.Q(p[30]));

	SEDFFX1 p_reg_31(
		.SI(p[25]),
		.SE(scan_en),
		.D(mpy_result[31]),
		.CK(clk),
		.E(n_6812),
		.Q(p[31]));

	SDFFRHQX1 pc_acc_reg(
		.SI(dp),
		.SE(scan_en),
		.D(n_3964),
		.CK(clk),
		.RN(n_7035),
		.Q(pc_acc));

	MXI2X1 i_4360(
		.S0(n_1439),
		.B(n_1114),
		.A(n_4222),
		.Y(n_3964));

	SDFFHQX1 null_op_reg(
		.SI(alu_cmd[2]),
		.SE(scan_en),
		.D(n_3973),
		.CK(clk),
		.Q(Q175));

	AND2X1 i_4369(
		.A(n_1109),
		.B(Q175),
		.Y(n_3973));

	SDFFHQX1 ar1_reg_0(
		.SI(Q175),
		.SE(scan_en),
		.D(n_4098),
		.CK(clk),
		.Q(ar1[0]));

	AOI21X1 i_4374(
		.A0(\nbus_424[0] ),
		.A1(ar1[0]),
		.B0(n_3978),
		.Y(n_3976));

	AOI21X1 i_4375(
		.A0(n_1061),
		.A1(n_781),
		.B0(\nbus_424[0] ),
		.Y(n_3978));

	SEDFFX1 ar1_reg_1(
		.SI(ar0[2]),
		.SE(scan_en),
		.D(\nbus_425[1] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[1]));

	SEDFFX1 ar1_reg_2(
		.SI(ar0[4]),
		.SE(scan_en),
		.D(\nbus_425[2] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[2]));

	SEDFFX1 ar1_reg_3(
		.SI(SPCASCAN_N29_present_state_1_),
		.SE(scan_en),
		.D(\nbus_425[3] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[3]));

	SEDFFX1 ar1_reg_4(
		.SI(ar0[5]),
		.SE(scan_en),
		.D(\nbus_425[4] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[4]));

	NAND2X1 i_2(
		.A(branch_stall),
		.B(phi_1),
		.Y(n_1103));

	SEDFFX1 ar1_reg_5(
		.SI(FE_PT3_),
		.SE(scan_en),
		.D(\nbus_425[5] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[5]));

	NOR3BX1 i_3521(
		.AN(n_1105),
		.B(n_859),
		.C(ir[3]),
		.Y(n_1104));

	SEDFFX1 ar1_reg_6(
		.SI(ar0[7]),
		.SE(scan_en),
		.D(\nbus_425[6] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[6]));

	NAND2BX1 i_2925(
		.AN(update_stall),
		.B(phi_5),
		.Y(n_1105));

	SEDFFX1 ar1_reg_7(
		.SI(ar0[6]),
		.SE(scan_en),
		.D(\nbus_425[7] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[7]));

	NOR2X1 i_2471(
		.A(n_832),
		.B(n_830),
		.Y(n_1106));

	SEDFFX1 ar1_reg_8(
		.SI(decode[13]),
		.SE(scan_en),
		.D(\nbus_425[8] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[8]));

	NAND4X1 i_3748(
		.A(phi_6),
		.B(n_7218),
		.C(n_429),
		.D(n_871),
		.Y(n_1107));

	SEDFFX1 ar1_reg_9(
		.SI(ar0[10]),
		.SE(scan_en),
		.D(\nbus_425[9] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[9]));

	AOI211X1 i_4043(
		.A0(n_1112),
		.A1(n_450),
		.B0(branch_stall_delay),
		.C0(branch_stall),
		.Y(n_1108));

	SEDFFX1 ar1_reg_10(
		.SI(ir[2]),
		.SE(scan_en),
		.D(\nbus_425[10] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[10]));

	OAI31X1 i_2860(
		.A0(n_717),
		.A1(n_1081),
		.A2(n_712),
		.B0(n_4076),
		.Y(n_1109));

	SEDFFX1 ar1_reg_11(
		.SI(ar0[11]),
		.SE(scan_en),
		.D(\nbus_425[11] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[11]));

	SEDFFX1 ar1_reg_12(
		.SI(ar0[8]),
		.SE(scan_en),
		.D(\nbus_425[12] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[12]));

	NAND2BX1 i_2475(
		.AN(n_813),
		.B(n_831),
		.Y(n_1111));

	SEDFFX1 ar1_reg_13(
		.SI(ar1[14]),
		.SE(scan_en),
		.D(\nbus_425[13] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[13]));

	NAND3BX1 i_2254(
		.AN(ir[2]),
		.B(ir[0]),
		.C(n_869),
		.Y(n_1112));

	SEDFFX1 ar1_reg_14(
		.SI(ar0[14]),
		.SE(scan_en),
		.D(\nbus_425[14] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[14]));

	SEDFFX1 ar1_reg_15(
		.SI(SPCASCAN_N28_read),
		.SE(scan_en),
		.D(\nbus_425[15] ),
		.CK(clk),
		.E(n_4099),
		.Q(ar1[15]));

	NAND2BX1 i_2698(
		.AN(n_793),
		.B(n_784),
		.Y(n_1114));

	INVX1 i_5175(
		.A(n_1001),
		.Y(n_4072));

	INVX1 i_5176(
		.A(n_998),
		.Y(n_4073));

	INVX1 i_5177(
		.A(n_995),
		.Y(n_4074));

	INVX1 i_5178(
		.A(n_1026),
		.Y(n_4075));

	INVX1 i_5179(
		.A(n_922),
		.Y(n_4076));

	INVX1 i_5180(
		.A(n_796),
		.Y(n_4077));

	INVX1 i_5181(
		.A(n_820),
		.Y(n_4078));

	INVX1 i_5182(
		.A(n_800),
		.Y(n_4079));

	INVX1 i_5183(
		.A(n_801),
		.Y(n_4080));

	INVX1 i_5184(
		.A(n_1111),
		.Y(n_4081));

	INVX1 i_5185(
		.A(n_804),
		.Y(n_4082));

	INVX1 i_5186(
		.A(n_1103),
		.Y(n_4083));

	INVX1 i_5187(
		.A(n_790),
		.Y(n_4084));

	INVX1 i_5188(
		.A(n_840),
		.Y(n_4085));

	INVX1 i_5189(
		.A(n_872),
		.Y(n_4086));

	INVX1 i_5190(
		.A(n_806),
		.Y(n_4087));

	INVX1 i_5191(
		.A(n_816),
		.Y(n_4088));

	INVX1 i_5192(
		.A(n_830),
		.Y(n_4089));

	INVX1 i_5193(
		.A(n_784),
		.Y(n_4090));

	INVX1 i_5194(
		.A(n_470),
		.Y(n_4091));

	INVX1 i_5195(
		.A(SPCASCAN_N32_two_cycle),
		.Y(n_4092));

	INVX1 i_5196(
		.A(n_3128),
		.Y(n_4093));

	INVX1 i_5197(
		.A(n_7384),
		.Y(n_4094));

	INVX1 i_5198(
		.A(n_3742),
		.Y(n_4095));

	INVX1 i_5199(
		.A(n_3748),
		.Y(n_4096));

	INVX1 i_5200(
		.A(\nbus_428[0] ),
		.Y(n_4097));

	INVX1 i_5201(
		.A(n_3976),
		.Y(n_4098));

	INVX1 i_5202(
		.A(\nbus_424[0] ),
		.Y(n_4099));

	INVX1 i_5203(
		.A(ir[8]),
		.Y(n_4100));

	INVX1 i_5204(
		.A(pc[12]),
		.Y(n_4101));

	INVX1 i_5205(
		.A(phi_1),
		.Y(n_4220));

	INVX1 i_5206(
		.A(reset),
		.Y(n_4221));

	INVX1 i_5207(
		.A(pc_acc),
		.Y(n_4222));

	INVX1 i_5208(
		.A(ovm),
		.Y(n_4223));

endmodule
module m16x16(
		a,
		b,
		y);

	input [15:0] a;
	input [15:0] b;
	output [31:0] y;




	AOI21X1 i_561(
		.A0(n_465),
		.A1(n_447),
		.B0(n_1024),
		.Y(y[1]));

	NAND3X1 i_558(
		.A(b[15]),
		.B(a[15]),
		.C(n_899),
		.Y(n_960));

	NAND2X1 i_557(
		.A(n_898),
		.B(n_897),
		.Y(n_959));

	NAND2X1 i_556(
		.A(n_896),
		.B(n_893),
		.Y(n_958));

	NAND2X1 i_555(
		.A(n_887),
		.B(n_892),
		.Y(n_957));

	NAND2X1 i_554(
		.A(n_886),
		.B(n_879),
		.Y(n_956));

	NAND2X1 i_553(
		.A(n_869),
		.B(n_878),
		.Y(n_955));

	NAND2X1 i_552(
		.A(n_857),
		.B(n_868),
		.Y(n_954));

	NAND2X1 i_551(
		.A(n_843),
		.B(n_856),
		.Y(n_953));

	NAND2X1 i_550(
		.A(n_842),
		.B(n_827),
		.Y(n_952));

	NAND2X1 i_549(
		.A(n_809),
		.B(n_826),
		.Y(n_951));

	NAND2X1 i_548(
		.A(n_789),
		.B(n_808),
		.Y(n_950));

	NAND2X1 i_547(
		.A(n_767),
		.B(n_788),
		.Y(n_949));

	NAND2X1 i_546(
		.A(n_743),
		.B(n_766),
		.Y(n_948));

	NAND2X1 i_545(
		.A(n_717),
		.B(n_742),
		.Y(n_947));

	NAND2X1 i_544(
		.A(n_689),
		.B(n_716),
		.Y(n_946));

	NAND2X1 i_543(
		.A(n_686),
		.B(n_688),
		.Y(n_945));

	NAND2X1 i_542(
		.A(n_635),
		.B(n_660),
		.Y(n_944));

	NAND2X1 i_541(
		.A(n_611),
		.B(n_634),
		.Y(n_943));

	NAND2X1 i_540(
		.A(n_589),
		.B(n_610),
		.Y(n_942));

	NAND2X1 i_539(
		.A(n_569),
		.B(n_588),
		.Y(n_941));

	NAND2X1 i_538(
		.A(n_566),
		.B(n_568),
		.Y(n_940));

	NAND2X1 i_537(
		.A(n_535),
		.B(n_550),
		.Y(n_939));

	NAND2X1 i_536(
		.A(n_521),
		.B(n_534),
		.Y(n_938));

	NAND2X1 i_535(
		.A(n_518),
		.B(n_520),
		.Y(n_937));

	NAND2X1 i_534(
		.A(n_499),
		.B(n_508),
		.Y(n_936));

	NAND2X1 i_533(
		.A(n_496),
		.B(n_498),
		.Y(n_935));

	NAND2X1 i_532(
		.A(n_485),
		.B(n_490),
		.Y(n_934));

	NAND2X1 i_531(
		.A(n_482),
		.B(n_484),
		.Y(n_933));

	NAND3X1 i_530(
		.A(b[2]),
		.B(a[0]),
		.C(n_480),
		.Y(n_932));

	NOR2X1 i_529(
		.A(n_465),
		.B(n_447),
		.Y(n_1024));

	AOI21X1 i_527(
		.A0(b[15]),
		.A1(a[15]),
		.B0(n_899),
		.Y(n_929));

	NOR2X1 i_526(
		.A(n_898),
		.B(n_897),
		.Y(n_928));

	NOR2X1 i_525(
		.A(n_896),
		.B(n_893),
		.Y(n_927));

	NOR2X1 i_524(
		.A(n_887),
		.B(n_892),
		.Y(n_926));

	NOR2X1 i_523(
		.A(n_886),
		.B(n_879),
		.Y(n_925));

	NOR2X1 i_522(
		.A(n_869),
		.B(n_878),
		.Y(n_924));

	NOR2X1 i_521(
		.A(n_857),
		.B(n_868),
		.Y(n_923));

	NOR2X1 i_520(
		.A(n_843),
		.B(n_856),
		.Y(n_922));

	NOR2X1 i_519(
		.A(n_842),
		.B(n_827),
		.Y(n_921));

	NOR2X1 i_518(
		.A(n_809),
		.B(n_826),
		.Y(n_920));

	NOR2X1 i_517(
		.A(n_789),
		.B(n_808),
		.Y(n_919));

	NOR2X1 i_516(
		.A(n_767),
		.B(n_788),
		.Y(n_918));

	NOR2X1 i_515(
		.A(n_743),
		.B(n_766),
		.Y(n_917));

	NOR2X1 i_514(
		.A(n_717),
		.B(n_742),
		.Y(n_916));

	NOR2X1 i_513(
		.A(n_689),
		.B(n_716),
		.Y(n_915));

	NOR2X1 i_512(
		.A(n_686),
		.B(n_688),
		.Y(n_914));

	NOR2X1 i_511(
		.A(n_635),
		.B(n_660),
		.Y(n_913));

	NOR2X1 i_510(
		.A(n_611),
		.B(n_634),
		.Y(n_912));

	NOR2X1 i_509(
		.A(n_589),
		.B(n_610),
		.Y(n_911));

	NOR2X1 i_508(
		.A(n_569),
		.B(n_588),
		.Y(n_910));

	NOR2X1 i_507(
		.A(n_566),
		.B(n_568),
		.Y(n_909));

	NOR2X1 i_506(
		.A(n_535),
		.B(n_550),
		.Y(n_908));

	NOR2X1 i_505(
		.A(n_521),
		.B(n_534),
		.Y(n_907));

	NOR2X1 i_504(
		.A(n_518),
		.B(n_520),
		.Y(n_906));

	NOR2X1 i_503(
		.A(n_499),
		.B(n_508),
		.Y(n_905));

	NOR2X1 i_502(
		.A(n_496),
		.B(n_498),
		.Y(n_904));

	NOR2X1 i_501(
		.A(n_485),
		.B(n_490),
		.Y(n_903));

	NOR2X1 i_500(
		.A(n_482),
		.B(n_484),
		.Y(n_902));

	AOI21X1 i_499(
		.A0(b[2]),
		.A1(a[0]),
		.B0(n_480),
		.Y(n_901));

	AND2X1 i_287(
		.A(b[0]),
		.B(a[15]),
		.Y(n_479));

	AND2X1 i_286(
		.A(b[0]),
		.B(a[14]),
		.Y(n_478));

	AND2X1 i_285(
		.A(b[0]),
		.B(a[13]),
		.Y(n_477));

	AND2X1 i_284(
		.A(b[0]),
		.B(a[12]),
		.Y(n_476));

	AND2X1 i_283(
		.A(b[0]),
		.B(a[11]),
		.Y(n_475));

	AND2X1 i_282(
		.A(b[0]),
		.B(a[10]),
		.Y(n_474));

	AND2X1 i_281(
		.A(b[0]),
		.B(a[9]),
		.Y(n_473));

	AND2X1 i_280(
		.A(b[0]),
		.B(a[8]),
		.Y(n_472));

	AND2X1 i_279(
		.A(b[0]),
		.B(a[7]),
		.Y(n_471));

	AND2X1 i_278(
		.A(b[0]),
		.B(a[6]),
		.Y(n_470));

	AND2X1 i_277(
		.A(b[0]),
		.B(a[5]),
		.Y(n_469));

	AND2X1 i_276(
		.A(b[0]),
		.B(a[4]),
		.Y(n_468));

	AND2X1 i_275(
		.A(b[0]),
		.B(a[3]),
		.Y(n_467));

	AND2X1 i_274(
		.A(b[0]),
		.B(a[2]),
		.Y(n_466));

	NAND2X1 i_273(
		.A(b[0]),
		.B(a[1]),
		.Y(n_465));

	AND2X1 i_272(
		.A(b[0]),
		.B(a[0]),
		.Y(y[0]));

	AOI31X1 i_563(
		.A0(b[2]),
		.A1(a[0]),
		.A2(n_480),
		.B0(n_901),
		.Y(n_965));

	AND2X1 i_270(
		.A(b[1]),
		.B(a[15]),
		.Y(n_462));

	AND2X1 i_269(
		.A(b[1]),
		.B(a[14]),
		.Y(n_461));

	AND2X1 i_268(
		.A(b[1]),
		.B(a[13]),
		.Y(n_460));

	AND2X1 i_267(
		.A(b[1]),
		.B(a[12]),
		.Y(n_459));

	AND2X1 i_266(
		.A(b[1]),
		.B(a[11]),
		.Y(n_458));

	AND2X1 i_265(
		.A(b[1]),
		.B(a[10]),
		.Y(n_457));

	AND2X1 i_264(
		.A(b[1]),
		.B(a[9]),
		.Y(n_456));

	AND2X1 i_263(
		.A(b[1]),
		.B(a[8]),
		.Y(n_455));

	AND2X1 i_262(
		.A(b[1]),
		.B(a[7]),
		.Y(n_454));

	AND2X1 i_261(
		.A(b[1]),
		.B(a[6]),
		.Y(n_453));

	AND2X1 i_260(
		.A(b[1]),
		.B(a[5]),
		.Y(n_452));

	AND2X1 i_259(
		.A(b[1]),
		.B(a[4]),
		.Y(n_451));

	AND2X1 i_258(
		.A(b[1]),
		.B(a[3]),
		.Y(n_450));

	AND2X1 i_257(
		.A(b[1]),
		.B(a[2]),
		.Y(n_449));

	AND2X1 i_256(
		.A(b[1]),
		.B(a[1]),
		.Y(n_448));

	NAND2X1 i_255(
		.A(b[1]),
		.B(a[0]),
		.Y(n_447));

	AOI21X1 i_565(
		.A0(n_482),
		.A1(n_484),
		.B0(n_902),
		.Y(n_967));

	AND2X1 i_253(
		.A(b[2]),
		.B(a[15]),
		.Y(n_445));

	AND2X1 i_252(
		.A(b[2]),
		.B(a[14]),
		.Y(n_444));

	AND2X1 i_251(
		.A(b[2]),
		.B(a[13]),
		.Y(n_443));

	AND2X1 i_250(
		.A(b[2]),
		.B(a[12]),
		.Y(n_442));

	AND2X1 i_249(
		.A(b[2]),
		.B(a[11]),
		.Y(n_441));

	AND2X1 i_248(
		.A(b[2]),
		.B(a[10]),
		.Y(n_440));

	AND2X1 i_247(
		.A(b[2]),
		.B(a[9]),
		.Y(n_439));

	AND2X1 i_246(
		.A(b[2]),
		.B(a[8]),
		.Y(n_438));

	AND2X1 i_245(
		.A(b[2]),
		.B(a[7]),
		.Y(n_437));

	AND2X1 i_244(
		.A(b[2]),
		.B(a[6]),
		.Y(n_436));

	AND2X1 i_243(
		.A(b[2]),
		.B(a[5]),
		.Y(n_435));

	AND2X1 i_242(
		.A(b[2]),
		.B(a[4]),
		.Y(n_434));

	AND2X1 i_241(
		.A(b[2]),
		.B(a[3]),
		.Y(n_433));

	AND2X1 i_240(
		.A(b[2]),
		.B(a[2]),
		.Y(n_432));

	AND2X1 i_239(
		.A(b[2]),
		.B(a[1]),
		.Y(n_431));

	AOI21X1 i_567(
		.A0(n_485),
		.A1(n_490),
		.B0(n_903),
		.Y(n_969));

	AND2X1 i_236(
		.A(b[3]),
		.B(a[15]),
		.Y(n_428));

	AND2X1 i_235(
		.A(b[3]),
		.B(a[14]),
		.Y(n_427));

	AND2X1 i_234(
		.A(b[3]),
		.B(a[13]),
		.Y(n_426));

	AND2X1 i_233(
		.A(b[3]),
		.B(a[12]),
		.Y(n_425));

	AND2X1 i_232(
		.A(b[3]),
		.B(a[11]),
		.Y(n_424));

	AND2X1 i_231(
		.A(b[3]),
		.B(a[10]),
		.Y(n_423));

	AND2X1 i_230(
		.A(b[3]),
		.B(a[9]),
		.Y(n_422));

	AND2X1 i_229(
		.A(b[3]),
		.B(a[8]),
		.Y(n_421));

	AND2X1 i_228(
		.A(b[3]),
		.B(a[7]),
		.Y(n_420));

	AND2X1 i_227(
		.A(b[3]),
		.B(a[6]),
		.Y(n_419));

	AND2X1 i_226(
		.A(b[3]),
		.B(a[5]),
		.Y(n_418));

	AND2X1 i_225(
		.A(b[3]),
		.B(a[4]),
		.Y(n_417));

	AND2X1 i_224(
		.A(b[3]),
		.B(a[3]),
		.Y(n_416));

	AND2X1 i_223(
		.A(b[3]),
		.B(a[2]),
		.Y(n_415));

	AND2X1 i_222(
		.A(b[3]),
		.B(a[1]),
		.Y(n_414));

	AND2X1 i_221(
		.A(b[3]),
		.B(a[0]),
		.Y(n_413));

	AOI21X1 i_569(
		.A0(n_496),
		.A1(n_498),
		.B0(n_904),
		.Y(n_971));

	AND2X1 i_219(
		.A(b[4]),
		.B(a[15]),
		.Y(n_411));

	AND2X1 i_218(
		.A(b[4]),
		.B(a[14]),
		.Y(n_410));

	AND2X1 i_217(
		.A(b[4]),
		.B(a[13]),
		.Y(n_409));

	AND2X1 i_216(
		.A(b[4]),
		.B(a[12]),
		.Y(n_408));

	AND2X1 i_215(
		.A(b[4]),
		.B(a[11]),
		.Y(n_407));

	AND2X1 i_214(
		.A(b[4]),
		.B(a[10]),
		.Y(n_406));

	AND2X1 i_213(
		.A(b[4]),
		.B(a[9]),
		.Y(n_405));

	AND2X1 i_212(
		.A(b[4]),
		.B(a[8]),
		.Y(n_404));

	AND2X1 i_211(
		.A(b[4]),
		.B(a[7]),
		.Y(n_403));

	AND2X1 i_210(
		.A(b[4]),
		.B(a[6]),
		.Y(n_402));

	AND2X1 i_209(
		.A(b[4]),
		.B(a[5]),
		.Y(n_401));

	AND2X1 i_208(
		.A(b[4]),
		.B(a[4]),
		.Y(n_400));

	AND2X1 i_207(
		.A(b[4]),
		.B(a[3]),
		.Y(n_399));

	AND2X1 i_206(
		.A(b[4]),
		.B(a[2]),
		.Y(n_398));

	AND2X1 i_205(
		.A(b[4]),
		.B(a[1]),
		.Y(n_397));

	AND2X1 i_204(
		.A(b[4]),
		.B(a[0]),
		.Y(n_396));

	AOI21X1 i_571(
		.A0(n_499),
		.A1(n_508),
		.B0(n_905),
		.Y(n_973));

	AND2X1 i_202(
		.A(b[5]),
		.B(a[15]),
		.Y(n_394));

	AND2X1 i_201(
		.A(b[5]),
		.B(a[14]),
		.Y(n_393));

	AND2X1 i_200(
		.A(b[5]),
		.B(a[13]),
		.Y(n_392));

	AND2X1 i_199(
		.A(b[5]),
		.B(a[12]),
		.Y(n_391));

	AND2X1 i_198(
		.A(b[5]),
		.B(a[11]),
		.Y(n_390));

	AND2X1 i_197(
		.A(b[5]),
		.B(a[10]),
		.Y(n_389));

	AND2X1 i_196(
		.A(b[5]),
		.B(a[9]),
		.Y(n_388));

	AND2X1 i_195(
		.A(b[5]),
		.B(a[8]),
		.Y(n_387));

	AND2X1 i_194(
		.A(b[5]),
		.B(a[7]),
		.Y(n_386));

	AND2X1 i_193(
		.A(b[5]),
		.B(a[6]),
		.Y(n_385));

	AND2X1 i_192(
		.A(b[5]),
		.B(a[5]),
		.Y(n_384));

	AND2X1 i_191(
		.A(b[5]),
		.B(a[4]),
		.Y(n_383));

	AND2X1 i_190(
		.A(b[5]),
		.B(a[3]),
		.Y(n_382));

	AND2X1 i_189(
		.A(b[5]),
		.B(a[2]),
		.Y(n_381));

	AND2X1 i_188(
		.A(b[5]),
		.B(a[1]),
		.Y(n_380));

	AND2X1 i_187(
		.A(b[5]),
		.B(a[0]),
		.Y(n_379));

	AOI21X1 i_573(
		.A0(n_518),
		.A1(n_520),
		.B0(n_906),
		.Y(n_975));

	AND2X1 i_185(
		.A(b[6]),
		.B(a[15]),
		.Y(n_377));

	AND2X1 i_184(
		.A(b[6]),
		.B(a[14]),
		.Y(n_376));

	AND2X1 i_183(
		.A(b[6]),
		.B(a[13]),
		.Y(n_375));

	AND2X1 i_182(
		.A(b[6]),
		.B(a[12]),
		.Y(n_374));

	AND2X1 i_181(
		.A(b[6]),
		.B(a[11]),
		.Y(n_373));

	AND2X1 i_180(
		.A(b[6]),
		.B(a[10]),
		.Y(n_372));

	AND2X1 i_179(
		.A(b[6]),
		.B(a[9]),
		.Y(n_371));

	AND2X1 i_178(
		.A(b[6]),
		.B(a[8]),
		.Y(n_370));

	AND2X1 i_177(
		.A(b[6]),
		.B(a[7]),
		.Y(n_369));

	AND2X1 i_176(
		.A(b[6]),
		.B(a[6]),
		.Y(n_368));

	AND2X1 i_175(
		.A(b[6]),
		.B(a[5]),
		.Y(n_367));

	AND2X1 i_174(
		.A(b[6]),
		.B(a[4]),
		.Y(n_366));

	AND2X1 i_173(
		.A(b[6]),
		.B(a[3]),
		.Y(n_365));

	AND2X1 i_172(
		.A(b[6]),
		.B(a[2]),
		.Y(n_364));

	AND2X1 i_171(
		.A(b[6]),
		.B(a[1]),
		.Y(n_363));

	AND2X1 i_170(
		.A(b[6]),
		.B(a[0]),
		.Y(n_362));

	AOI21X1 i_575(
		.A0(n_521),
		.A1(n_534),
		.B0(n_907),
		.Y(n_977));

	AND2X1 i_168(
		.A(b[7]),
		.B(a[15]),
		.Y(n_360));

	AND2X1 i_167(
		.A(b[7]),
		.B(a[14]),
		.Y(n_359));

	AND2X1 i_166(
		.A(b[7]),
		.B(a[13]),
		.Y(n_358));

	AND2X1 i_165(
		.A(b[7]),
		.B(a[12]),
		.Y(n_357));

	AND2X1 i_164(
		.A(b[7]),
		.B(a[11]),
		.Y(n_356));

	AND2X1 i_163(
		.A(b[7]),
		.B(a[10]),
		.Y(n_355));

	AND2X1 i_162(
		.A(b[7]),
		.B(a[9]),
		.Y(n_354));

	AND2X1 i_161(
		.A(b[7]),
		.B(a[8]),
		.Y(n_353));

	AND2X1 i_160(
		.A(b[7]),
		.B(a[7]),
		.Y(n_352));

	AND2X1 i_159(
		.A(b[7]),
		.B(a[6]),
		.Y(n_351));

	AND2X1 i_158(
		.A(b[7]),
		.B(a[5]),
		.Y(n_350));

	AND2X1 i_157(
		.A(b[7]),
		.B(a[4]),
		.Y(n_349));

	AND2X1 i_156(
		.A(b[7]),
		.B(a[3]),
		.Y(n_348));

	AND2X1 i_155(
		.A(b[7]),
		.B(a[2]),
		.Y(n_347));

	AND2X1 i_154(
		.A(b[7]),
		.B(a[1]),
		.Y(n_346));

	AND2X1 i_153(
		.A(b[7]),
		.B(a[0]),
		.Y(n_345));

	AOI21X1 i_577(
		.A0(n_535),
		.A1(n_550),
		.B0(n_908),
		.Y(n_979));

	AND2X1 i_151(
		.A(b[8]),
		.B(a[15]),
		.Y(n_343));

	AND2X1 i_150(
		.A(b[8]),
		.B(a[14]),
		.Y(n_342));

	AND2X1 i_149(
		.A(b[8]),
		.B(a[13]),
		.Y(n_341));

	AND2X1 i_148(
		.A(b[8]),
		.B(a[12]),
		.Y(n_340));

	AND2X1 i_147(
		.A(b[8]),
		.B(a[11]),
		.Y(n_339));

	AND2X1 i_146(
		.A(b[8]),
		.B(a[10]),
		.Y(n_338));

	AND2X1 i_145(
		.A(b[8]),
		.B(a[9]),
		.Y(n_337));

	AND2X1 i_144(
		.A(b[8]),
		.B(a[8]),
		.Y(n_336));

	AND2X1 i_143(
		.A(b[8]),
		.B(a[7]),
		.Y(n_335));

	AND2X1 i_142(
		.A(b[8]),
		.B(a[6]),
		.Y(n_334));

	AND2X1 i_141(
		.A(b[8]),
		.B(a[5]),
		.Y(n_333));

	AND2X1 i_140(
		.A(b[8]),
		.B(a[4]),
		.Y(n_332));

	AND2X1 i_139(
		.A(b[8]),
		.B(a[3]),
		.Y(n_331));

	AND2X1 i_138(
		.A(b[8]),
		.B(a[2]),
		.Y(n_330));

	AND2X1 i_137(
		.A(b[8]),
		.B(a[1]),
		.Y(n_329));

	AND2X1 i_136(
		.A(b[8]),
		.B(a[0]),
		.Y(n_328));

	AOI21X1 i_579(
		.A0(n_566),
		.A1(n_568),
		.B0(n_909),
		.Y(n_981));

	AND2X1 i_134(
		.A(b[9]),
		.B(a[15]),
		.Y(n_326));

	AND2X1 i_133(
		.A(b[9]),
		.B(a[14]),
		.Y(n_325));

	AND2X1 i_132(
		.A(b[9]),
		.B(a[13]),
		.Y(n_324));

	AND2X1 i_131(
		.A(b[9]),
		.B(a[12]),
		.Y(n_323));

	AND2X1 i_130(
		.A(b[9]),
		.B(a[11]),
		.Y(n_322));

	AND2X1 i_129(
		.A(b[9]),
		.B(a[10]),
		.Y(n_321));

	AND2X1 i_128(
		.A(b[9]),
		.B(a[9]),
		.Y(n_320));

	AND2X1 i_127(
		.A(b[9]),
		.B(a[8]),
		.Y(n_319));

	AND2X1 i_126(
		.A(b[9]),
		.B(a[7]),
		.Y(n_318));

	AND2X1 i_125(
		.A(b[9]),
		.B(a[6]),
		.Y(n_317));

	AND2X1 i_124(
		.A(b[9]),
		.B(a[5]),
		.Y(n_316));

	AND2X1 i_123(
		.A(b[9]),
		.B(a[4]),
		.Y(n_315));

	AND2X1 i_122(
		.A(b[9]),
		.B(a[3]),
		.Y(n_314));

	AND2X1 i_121(
		.A(b[9]),
		.B(a[2]),
		.Y(n_313));

	AND2X1 i_120(
		.A(b[9]),
		.B(a[1]),
		.Y(n_312));

	AND2X1 i_119(
		.A(b[9]),
		.B(a[0]),
		.Y(n_311));

	AOI21X1 i_581(
		.A0(n_569),
		.A1(n_588),
		.B0(n_910),
		.Y(n_983));

	AND2X1 i_117(
		.A(b[10]),
		.B(a[15]),
		.Y(n_309));

	AND2X1 i_116(
		.A(b[10]),
		.B(a[14]),
		.Y(n_308));

	AND2X1 i_115(
		.A(b[10]),
		.B(a[13]),
		.Y(n_307));

	AND2X1 i_114(
		.A(b[10]),
		.B(a[12]),
		.Y(n_306));

	AND2X1 i_113(
		.A(b[10]),
		.B(a[11]),
		.Y(n_305));

	AND2X1 i_112(
		.A(b[10]),
		.B(a[10]),
		.Y(n_304));

	AND2X1 i_111(
		.A(b[10]),
		.B(a[9]),
		.Y(n_303));

	AND2X1 i_110(
		.A(b[10]),
		.B(a[8]),
		.Y(n_302));

	AND2X1 i_109(
		.A(b[10]),
		.B(a[7]),
		.Y(n_301));

	AND2X1 i_108(
		.A(b[10]),
		.B(a[6]),
		.Y(n_300));

	AND2X1 i_107(
		.A(b[10]),
		.B(a[5]),
		.Y(n_299));

	AND2X1 i_106(
		.A(b[10]),
		.B(a[4]),
		.Y(n_298));

	AND2X1 i_105(
		.A(b[10]),
		.B(a[3]),
		.Y(n_297));

	AND2X1 i_104(
		.A(b[10]),
		.B(a[2]),
		.Y(n_296));

	AND2X1 i_103(
		.A(b[10]),
		.B(a[1]),
		.Y(n_295));

	AND2X1 i_102(
		.A(b[10]),
		.B(a[0]),
		.Y(n_294));

	AOI21X1 i_583(
		.A0(n_589),
		.A1(n_610),
		.B0(n_911),
		.Y(n_985));

	AND2X1 i_100(
		.A(b[11]),
		.B(a[15]),
		.Y(n_292));

	AND2X1 i_99(
		.A(b[11]),
		.B(a[14]),
		.Y(n_291));

	AND2X1 i_98(
		.A(b[11]),
		.B(a[13]),
		.Y(n_290));

	AND2X1 i_97(
		.A(b[11]),
		.B(a[12]),
		.Y(n_289));

	AND2X1 i_96(
		.A(b[11]),
		.B(a[11]),
		.Y(n_288));

	AND2X1 i_95(
		.A(b[11]),
		.B(a[10]),
		.Y(n_287));

	AND2X1 i_94(
		.A(b[11]),
		.B(a[9]),
		.Y(n_286));

	AND2X1 i_93(
		.A(b[11]),
		.B(a[8]),
		.Y(n_285));

	AND2X1 i_92(
		.A(b[11]),
		.B(a[7]),
		.Y(n_284));

	AND2X1 i_91(
		.A(b[11]),
		.B(a[6]),
		.Y(n_283));

	AND2X1 i_90(
		.A(b[11]),
		.B(a[5]),
		.Y(n_282));

	AND2X1 i_89(
		.A(b[11]),
		.B(a[4]),
		.Y(n_281));

	AND2X1 i_88(
		.A(b[11]),
		.B(a[3]),
		.Y(n_280));

	AND2X1 i_87(
		.A(b[11]),
		.B(a[2]),
		.Y(n_279));

	AND2X1 i_86(
		.A(b[11]),
		.B(a[1]),
		.Y(n_278));

	AND2X1 i_85(
		.A(b[11]),
		.B(a[0]),
		.Y(n_277));

	AOI21X1 i_585(
		.A0(n_611),
		.A1(n_634),
		.B0(n_912),
		.Y(n_987));

	AND2X1 i_83(
		.A(b[12]),
		.B(a[15]),
		.Y(n_275));

	AND2X1 i_82(
		.A(b[12]),
		.B(a[14]),
		.Y(n_274));

	AND2X1 i_81(
		.A(b[12]),
		.B(a[13]),
		.Y(n_273));

	AND2X1 i_80(
		.A(b[12]),
		.B(a[12]),
		.Y(n_272));

	AND2X1 i_79(
		.A(b[12]),
		.B(a[11]),
		.Y(n_271));

	AND2X1 i_78(
		.A(b[12]),
		.B(a[10]),
		.Y(n_270));

	AND2X1 i_77(
		.A(b[12]),
		.B(a[9]),
		.Y(n_269));

	AND2X1 i_76(
		.A(b[12]),
		.B(a[8]),
		.Y(n_268));

	AND2X1 i_75(
		.A(b[12]),
		.B(a[7]),
		.Y(n_267));

	AND2X1 i_74(
		.A(b[12]),
		.B(a[6]),
		.Y(n_266));

	AND2X1 i_73(
		.A(b[12]),
		.B(a[5]),
		.Y(n_265));

	AND2X1 i_72(
		.A(b[12]),
		.B(a[4]),
		.Y(n_264));

	AND2X1 i_71(
		.A(b[12]),
		.B(a[3]),
		.Y(n_263));

	AND2X1 i_70(
		.A(b[12]),
		.B(a[2]),
		.Y(n_262));

	AND2X1 i_69(
		.A(b[12]),
		.B(a[1]),
		.Y(n_261));

	AND2X1 i_68(
		.A(b[12]),
		.B(a[0]),
		.Y(n_260));

	AOI21X1 i_587(
		.A0(n_635),
		.A1(n_660),
		.B0(n_913),
		.Y(n_989));

	AND2X1 i_66(
		.A(b[13]),
		.B(a[15]),
		.Y(n_258));

	AND2X1 i_65(
		.A(b[13]),
		.B(a[14]),
		.Y(n_257));

	AND2X1 i_64(
		.A(b[13]),
		.B(a[13]),
		.Y(n_256));

	AND2X1 i_63(
		.A(b[13]),
		.B(a[12]),
		.Y(n_255));

	AND2X1 i_62(
		.A(b[13]),
		.B(a[11]),
		.Y(n_254));

	AND2X1 i_61(
		.A(b[13]),
		.B(a[10]),
		.Y(n_253));

	AND2X1 i_60(
		.A(b[13]),
		.B(a[9]),
		.Y(n_252));

	AND2X1 i_59(
		.A(b[13]),
		.B(a[8]),
		.Y(n_251));

	AND2X1 i_58(
		.A(b[13]),
		.B(a[7]),
		.Y(n_250));

	AND2X1 i_57(
		.A(b[13]),
		.B(a[6]),
		.Y(n_249));

	AND2X1 i_56(
		.A(b[13]),
		.B(a[5]),
		.Y(n_248));

	AND2X1 i_55(
		.A(b[13]),
		.B(a[4]),
		.Y(n_247));

	AND2X1 i_54(
		.A(b[13]),
		.B(a[3]),
		.Y(n_246));

	AND2X1 i_53(
		.A(b[13]),
		.B(a[2]),
		.Y(n_245));

	AND2X1 i_52(
		.A(b[13]),
		.B(a[1]),
		.Y(n_244));

	AND2X1 i_51(
		.A(b[13]),
		.B(a[0]),
		.Y(n_243));

	AOI21X1 i_589(
		.A0(n_686),
		.A1(n_688),
		.B0(n_914),
		.Y(n_991));

	AND2X1 i_49(
		.A(b[14]),
		.B(a[15]),
		.Y(n_241));

	AND2X1 i_48(
		.A(b[14]),
		.B(a[14]),
		.Y(n_240));

	AND2X1 i_47(
		.A(b[14]),
		.B(a[13]),
		.Y(n_239));

	AND2X1 i_46(
		.A(b[14]),
		.B(a[12]),
		.Y(n_238));

	AND2X1 i_45(
		.A(b[14]),
		.B(a[11]),
		.Y(n_237));

	AND2X1 i_44(
		.A(b[14]),
		.B(a[10]),
		.Y(n_236));

	AND2X1 i_43(
		.A(b[14]),
		.B(a[9]),
		.Y(n_235));

	AND2X1 i_42(
		.A(b[14]),
		.B(a[8]),
		.Y(n_234));

	AND2X1 i_41(
		.A(b[14]),
		.B(a[7]),
		.Y(n_233));

	AND2X1 i_40(
		.A(b[14]),
		.B(a[6]),
		.Y(n_232));

	AND2X1 i_39(
		.A(b[14]),
		.B(a[5]),
		.Y(n_231));

	AND2X1 i_38(
		.A(b[14]),
		.B(a[4]),
		.Y(n_230));

	AND2X1 i_37(
		.A(b[14]),
		.B(a[3]),
		.Y(n_229));

	AND2X1 i_36(
		.A(b[14]),
		.B(a[2]),
		.Y(n_228));

	AND2X1 i_35(
		.A(b[14]),
		.B(a[1]),
		.Y(n_227));

	AND2X1 i_34(
		.A(b[14]),
		.B(a[0]),
		.Y(n_226));

	AOI21X1 i_591(
		.A0(n_689),
		.A1(n_716),
		.B0(n_915),
		.Y(n_993));

	AND2X1 i_31(
		.A(b[15]),
		.B(a[14]),
		.Y(n_223));

	AND2X1 i_30(
		.A(b[15]),
		.B(a[13]),
		.Y(n_222));

	AND2X1 i_29(
		.A(b[15]),
		.B(a[12]),
		.Y(n_221));

	AND2X1 i_28(
		.A(b[15]),
		.B(a[11]),
		.Y(n_220));

	AND2X1 i_27(
		.A(b[15]),
		.B(a[10]),
		.Y(n_219));

	AND2X1 i_26(
		.A(b[15]),
		.B(a[9]),
		.Y(n_218));

	AND2X1 i_25(
		.A(b[15]),
		.B(a[8]),
		.Y(n_217));

	AND2X1 i_24(
		.A(b[15]),
		.B(a[7]),
		.Y(n_216));

	AND2X1 i_23(
		.A(b[15]),
		.B(a[6]),
		.Y(n_215));

	AND2X1 i_22(
		.A(b[15]),
		.B(a[5]),
		.Y(n_214));

	AND2X1 i_21(
		.A(b[15]),
		.B(a[4]),
		.Y(n_213));

	AND2X1 i_20(
		.A(b[15]),
		.B(a[3]),
		.Y(n_212));

	AND2X1 i_19(
		.A(b[15]),
		.B(a[2]),
		.Y(n_211));

	AND2X1 i_18(
		.A(b[15]),
		.B(a[1]),
		.Y(n_210));

	AND2X1 i_17(
		.A(b[15]),
		.B(a[0]),
		.Y(n_209));

	AOI21X1 i_593(
		.A0(n_717),
		.A1(n_742),
		.B0(n_916),
		.Y(n_995));

	AOI21X1 i_595(
		.A0(n_743),
		.A1(n_766),
		.B0(n_917),
		.Y(n_997));

	AOI21X1 i_597(
		.A0(n_767),
		.A1(n_788),
		.B0(n_918),
		.Y(n_999));

	AOI21X1 i_599(
		.A0(n_789),
		.A1(n_808),
		.B0(n_919),
		.Y(n_1001));

	AOI21X1 i_601(
		.A0(n_809),
		.A1(n_826),
		.B0(n_920),
		.Y(n_1003));

	AOI21X1 i_603(
		.A0(n_842),
		.A1(n_827),
		.B0(n_921),
		.Y(n_1005));

	AOI21X1 i_605(
		.A0(n_843),
		.A1(n_856),
		.B0(n_922),
		.Y(n_1007));

	AOI21X1 i_607(
		.A0(n_857),
		.A1(n_868),
		.B0(n_923),
		.Y(n_1009));

	AOI21X1 i_609(
		.A0(n_869),
		.A1(n_878),
		.B0(n_924),
		.Y(n_1011));

	AOI21X1 i_611(
		.A0(n_886),
		.A1(n_879),
		.B0(n_925),
		.Y(n_1013));

	AOI21X1 i_613(
		.A0(n_887),
		.A1(n_892),
		.B0(n_926),
		.Y(n_1015));

	AOI21X1 i_615(
		.A0(n_896),
		.A1(n_893),
		.B0(n_927),
		.Y(n_1017));

	AOI21X1 i_617(
		.A0(n_898),
		.A1(n_897),
		.B0(n_928),
		.Y(n_1019));

	AOI31X1 i_619(
		.A0(b[15]),
		.A1(a[15]),
		.A2(n_899),
		.B0(n_929),
		.Y(n_1021));

	NOR2X1 i_654(
		.A(n_902),
		.B(n_901),
		.Y(n_1056));

	NOR2X1 i_655(
		.A(n_903),
		.B(n_902),
		.Y(n_1057));

	NOR2X1 i_656(
		.A(n_904),
		.B(n_903),
		.Y(n_1058));

	XNOR2X1 i_893(
		.A(n_965),
		.B(n_931),
		.Y(y[2]));

	NOR2X1 i_657(
		.A(n_905),
		.B(n_904),
		.Y(n_1059));

	NOR2X1 i_658(
		.A(n_906),
		.B(n_905),
		.Y(n_1060));

	NOR2X1 i_659(
		.A(n_907),
		.B(n_906),
		.Y(n_1061));

	AOI21X1 i_894(
		.A0(n_967),
		.A1(n_1025),
		.B0(n_5393),
		.Y(y[3]));

	NOR2X1 i_6310(
		.A(n_967),
		.B(n_1025),
		.Y(n_5393));

	NOR2X1 i_660(
		.A(n_908),
		.B(n_907),
		.Y(n_1062));

	NOR2X1 i_661(
		.A(n_909),
		.B(n_908),
		.Y(n_1063));

	NOR2X1 i_662(
		.A(n_910),
		.B(n_909),
		.Y(n_1064));

	XNOR2X1 i_895(
		.A(n_969),
		.B(n_1086),
		.Y(y[4]));

	NOR2X1 i_663(
		.A(n_911),
		.B(n_910),
		.Y(n_1065));

	NOR2X1 i_664(
		.A(n_912),
		.B(n_911),
		.Y(n_1066));

	NOR2X1 i_665(
		.A(n_913),
		.B(n_912),
		.Y(n_1067));

	XNOR2X1 i_896(
		.A(n_971),
		.B(n_1087),
		.Y(y[5]));

	NOR2X1 i_666(
		.A(n_914),
		.B(n_913),
		.Y(n_1068));

	NOR2X1 i_667(
		.A(n_915),
		.B(n_914),
		.Y(n_1069));

	NOR2X1 i_668(
		.A(n_916),
		.B(n_915),
		.Y(n_1070));

	AOI21X1 i_897(
		.A0(n_973),
		.A1(n_1148),
		.B0(n_5408),
		.Y(y[6]));

	NOR2X1 i_6325(
		.A(n_973),
		.B(n_1148),
		.Y(n_5408));

	NOR2X1 i_669(
		.A(n_917),
		.B(n_916),
		.Y(n_1071));

	NOR2X1 i_670(
		.A(n_918),
		.B(n_917),
		.Y(n_1072));

	NOR2X1 i_671(
		.A(n_919),
		.B(n_918),
		.Y(n_1073));

	AOI21X1 i_898(
		.A0(n_975),
		.A1(n_1149),
		.B0(n_5413),
		.Y(y[7]));

	NOR2X1 i_6330(
		.A(n_975),
		.B(n_1149),
		.Y(n_5413));

	NOR2X1 i_672(
		.A(n_920),
		.B(n_919),
		.Y(n_1074));

	NOR2X1 i_673(
		.A(n_921),
		.B(n_920),
		.Y(n_1075));

	NOR2X1 i_674(
		.A(n_922),
		.B(n_921),
		.Y(n_1076));

	AOI21X1 i_899(
		.A0(n_977),
		.A1(n_1150),
		.B0(n_5418),
		.Y(y[8]));

	NOR2X1 i_6335(
		.A(n_977),
		.B(n_1150),
		.Y(n_5418));

	NOR2X1 i_675(
		.A(n_923),
		.B(n_922),
		.Y(n_1077));

	NOR2X1 i_676(
		.A(n_924),
		.B(n_923),
		.Y(n_1078));

	NOR2X1 i_677(
		.A(n_925),
		.B(n_924),
		.Y(n_1079));

	AOI21X1 i_900(
		.A0(n_979),
		.A1(n_1151),
		.B0(n_5423),
		.Y(y[9]));

	NOR2X1 i_6340(
		.A(n_979),
		.B(n_1151),
		.Y(n_5423));

	NOR2X1 i_678(
		.A(n_926),
		.B(n_925),
		.Y(n_1080));

	NOR2X1 i_679(
		.A(n_927),
		.B(n_926),
		.Y(n_1081));

	NOR2X1 i_680(
		.A(n_928),
		.B(n_927),
		.Y(n_1082));

	XNOR2X1 i_901(
		.A(n_981),
		.B(n_1212),
		.Y(y[10]));

	NOR2X1 i_681(
		.A(n_929),
		.B(n_928),
		.Y(n_1083));

	NAND2X1 i_716(
		.A(n_1058),
		.B(n_1056),
		.Y(n_1118));

	NAND2X1 i_717(
		.A(n_1059),
		.B(n_1057),
		.Y(n_1119));

	XNOR2X1 i_902(
		.A(n_983),
		.B(n_1213),
		.Y(y[11]));

	NAND2X1 i_718(
		.A(n_1060),
		.B(n_1058),
		.Y(n_1120));

	NAND2X1 i_719(
		.A(n_1061),
		.B(n_1059),
		.Y(n_1121));

	NAND2X1 i_720(
		.A(n_1062),
		.B(n_1060),
		.Y(n_1122));

	XNOR2X1 i_903(
		.A(n_985),
		.B(n_1214),
		.Y(y[12]));

	NAND2X1 i_721(
		.A(n_1063),
		.B(n_1061),
		.Y(n_1123));

	NAND2X1 i_722(
		.A(n_1064),
		.B(n_1062),
		.Y(n_1124));

	NAND2X1 i_723(
		.A(n_1065),
		.B(n_1063),
		.Y(n_1125));

	XNOR2X1 i_904(
		.A(n_987),
		.B(n_1215),
		.Y(y[13]));

	NAND2X1 i_724(
		.A(n_1066),
		.B(n_1064),
		.Y(n_1126));

	NAND2X1 i_725(
		.A(n_1067),
		.B(n_1065),
		.Y(n_1127));

	NAND2X1 i_726(
		.A(n_1068),
		.B(n_1066),
		.Y(n_1128));

	XNOR2X1 i_905(
		.A(n_989),
		.B(n_1216),
		.Y(y[14]));

	NAND2X1 i_727(
		.A(n_1069),
		.B(n_1067),
		.Y(n_1129));

	NAND2X1 i_728(
		.A(n_1070),
		.B(n_1068),
		.Y(n_1130));

	NAND2X1 i_729(
		.A(n_1071),
		.B(n_1069),
		.Y(n_1131));

	XNOR2X1 i_906(
		.A(n_991),
		.B(n_1217),
		.Y(y[15]));

	NAND2X1 i_730(
		.A(n_1072),
		.B(n_1070),
		.Y(n_1132));

	NAND2X1 i_731(
		.A(n_1073),
		.B(n_1071),
		.Y(n_1133));

	NAND2X1 i_732(
		.A(n_1074),
		.B(n_1072),
		.Y(n_1134));

	XNOR2X1 i_907(
		.A(n_993),
		.B(n_1218),
		.Y(y[16]));

	NAND2X1 i_733(
		.A(n_1075),
		.B(n_1073),
		.Y(n_1135));

	NAND2X1 i_734(
		.A(n_1076),
		.B(n_1074),
		.Y(n_1136));

	NAND2X1 i_735(
		.A(n_1077),
		.B(n_1075),
		.Y(n_1137));

	XNOR2X1 i_908(
		.A(n_995),
		.B(n_1219),
		.Y(y[17]));

	NAND2X1 i_736(
		.A(n_1078),
		.B(n_1076),
		.Y(n_1138));

	NAND2X1 i_737(
		.A(n_1079),
		.B(n_1077),
		.Y(n_1139));

	NAND2X1 i_738(
		.A(n_1080),
		.B(n_1078),
		.Y(n_1140));

	AOI21X1 i_909(
		.A0(n_997),
		.A1(n_1280),
		.B0(n_5468),
		.Y(y[18]));

	NOR2X1 i_6385(
		.A(n_997),
		.B(n_1280),
		.Y(n_5468));

	NAND2X1 i_739(
		.A(n_1081),
		.B(n_1079),
		.Y(n_1141));

	NAND2X1 i_740(
		.A(n_1082),
		.B(n_1080),
		.Y(n_1142));

	NAND2X1 i_741(
		.A(n_1083),
		.B(n_1081),
		.Y(n_1143));

	AOI21X1 i_910(
		.A0(n_999),
		.A1(n_1281),
		.B0(n_5473),
		.Y(y[19]));

	NOR2X1 i_6390(
		.A(n_999),
		.B(n_1281),
		.Y(n_5473));

	NOR2X1 i_780(
		.A(n_1122),
		.B(n_1118),
		.Y(n_1182));

	NOR2X1 i_781(
		.A(n_1123),
		.B(n_1119),
		.Y(n_1183));

	NOR2X1 i_782(
		.A(n_1124),
		.B(n_1120),
		.Y(n_1184));

	AOI21X1 i_911(
		.A0(n_1001),
		.A1(n_1282),
		.B0(n_5478),
		.Y(y[20]));

	NOR2X1 i_6395(
		.A(n_1001),
		.B(n_1282),
		.Y(n_5478));

	NOR2X1 i_783(
		.A(n_1125),
		.B(n_1121),
		.Y(n_1185));

	NOR2X1 i_784(
		.A(n_1126),
		.B(n_1122),
		.Y(n_1186));

	NOR2X1 i_785(
		.A(n_1127),
		.B(n_1123),
		.Y(n_1187));

	AOI21X1 i_912(
		.A0(n_1003),
		.A1(n_1283),
		.B0(n_5483),
		.Y(y[21]));

	NOR2X1 i_6400(
		.A(n_1003),
		.B(n_1283),
		.Y(n_5483));

	NOR2X1 i_786(
		.A(n_1128),
		.B(n_1124),
		.Y(n_1188));

	NOR2X1 i_787(
		.A(n_1129),
		.B(n_1125),
		.Y(n_1189));

	NOR2X1 i_788(
		.A(n_1130),
		.B(n_1126),
		.Y(n_1190));

	AOI21X1 i_913(
		.A0(n_1005),
		.A1(n_1284),
		.B0(n_5488),
		.Y(y[22]));

	NOR2X1 i_6405(
		.A(n_1005),
		.B(n_1284),
		.Y(n_5488));

	NOR2X1 i_789(
		.A(n_1131),
		.B(n_1127),
		.Y(n_1191));

	NOR2X1 i_790(
		.A(n_1132),
		.B(n_1128),
		.Y(n_1192));

	NOR2X1 i_791(
		.A(n_1133),
		.B(n_1129),
		.Y(n_1193));

	AOI21X1 i_914(
		.A0(n_1007),
		.A1(n_1285),
		.B0(n_5493),
		.Y(y[23]));

	NOR2X1 i_6410(
		.A(n_1007),
		.B(n_1285),
		.Y(n_5493));

	NOR2X1 i_792(
		.A(n_1134),
		.B(n_1130),
		.Y(n_1194));

	NOR2X1 i_793(
		.A(n_1135),
		.B(n_1131),
		.Y(n_1195));

	NOR2X1 i_794(
		.A(n_1136),
		.B(n_1132),
		.Y(n_1196));

	AOI21X1 i_915(
		.A0(n_1009),
		.A1(n_1286),
		.B0(n_5498),
		.Y(y[24]));

	NOR2X1 i_6415(
		.A(n_1009),
		.B(n_1286),
		.Y(n_5498));

	NOR2X1 i_795(
		.A(n_1137),
		.B(n_1133),
		.Y(n_1197));

	NOR2X1 i_796(
		.A(n_1138),
		.B(n_1134),
		.Y(n_1198));

	NOR2X1 i_797(
		.A(n_1139),
		.B(n_1135),
		.Y(n_1199));

	AOI21X1 i_916(
		.A0(n_1011),
		.A1(n_1287),
		.B0(n_5503),
		.Y(y[25]));

	NOR2X1 i_6420(
		.A(n_1011),
		.B(n_1287),
		.Y(n_5503));

	NOR2X1 i_798(
		.A(n_1140),
		.B(n_1136),
		.Y(n_1200));

	NOR2X1 i_799(
		.A(n_1141),
		.B(n_1137),
		.Y(n_1201));

	NOR2X1 i_800(
		.A(n_1142),
		.B(n_1138),
		.Y(n_1202));

	AOI21X1 i_917(
		.A0(n_1013),
		.A1(n_1288),
		.B0(n_5508),
		.Y(y[26]));

	NOR2X1 i_6425(
		.A(n_1013),
		.B(n_1288),
		.Y(n_5508));

	NOR2X1 i_801(
		.A(n_1143),
		.B(n_1139),
		.Y(n_1203));

	NAND2X1 i_848(
		.A(n_1182),
		.B(n_1190),
		.Y(n_1250));

	NAND2X1 i_849(
		.A(n_1183),
		.B(n_1191),
		.Y(n_1251));

	AOI21X1 i_918(
		.A0(n_1015),
		.A1(n_1289),
		.B0(n_5513),
		.Y(y[27]));

	NOR2X1 i_6430(
		.A(n_1015),
		.B(n_1289),
		.Y(n_5513));

	NAND2X1 i_850(
		.A(n_1184),
		.B(n_1192),
		.Y(n_1252));

	NAND2X1 i_851(
		.A(n_1185),
		.B(n_1193),
		.Y(n_1253));

	NAND2X1 i_852(
		.A(n_1186),
		.B(n_1194),
		.Y(n_1254));

	AOI21X1 i_919(
		.A0(n_1017),
		.A1(n_1290),
		.B0(n_5518),
		.Y(y[28]));

	NOR2X1 i_6435(
		.A(n_1017),
		.B(n_1290),
		.Y(n_5518));

	NAND2X1 i_853(
		.A(n_1195),
		.B(n_1187),
		.Y(n_1255));

	NAND2X1 i_854(
		.A(n_1188),
		.B(n_1196),
		.Y(n_1256));

	NAND2X1 i_855(
		.A(n_1189),
		.B(n_1197),
		.Y(n_1257));

	AOI21X1 i_920(
		.A0(n_1019),
		.A1(n_1291),
		.B0(n_5523),
		.Y(y[29]));

	NOR2X1 i_6440(
		.A(n_1019),
		.B(n_1291),
		.Y(n_5523));

	NAND2X1 i_856(
		.A(n_1190),
		.B(n_1198),
		.Y(n_1258));

	NAND2X1 i_857(
		.A(n_1191),
		.B(n_1199),
		.Y(n_1259));

	NAND4BXL i_858(
		.AN(n_1136),
		.B(n_1080),
		.C(n_1078),
		.D(n_1192),
		.Y(n_1260));

	AOI21X1 i_921(
		.A0(n_1021),
		.A1(n_1292),
		.B0(n_5528),
		.Y(y[30]));

	NOR2X1 i_6445(
		.A(n_1021),
		.B(n_1292),
		.Y(n_5528));

	NAND4BXL i_859(
		.AN(n_1137),
		.B(n_1081),
		.C(n_1079),
		.D(n_1193),
		.Y(n_1261));

	NAND4BXL i_860(
		.AN(n_1138),
		.B(n_1082),
		.C(n_1080),
		.D(n_1194),
		.Y(n_1262));

	NAND2X1 i_861(
		.A(n_1203),
		.B(n_1195),
		.Y(n_1263));

	INVX1 i_6930(
		.A(n_1151),
		.Y(n_1211));

	INVX1 i_6931(
		.A(n_1150),
		.Y(n_1210));

	INVX1 i_6932(
		.A(n_1149),
		.Y(n_1209));

	INVX1 i_6933(
		.A(n_1148),
		.Y(n_1208));

	INVX1 i_6934(
		.A(n_1025),
		.Y(n_1085));

	INVX1 i_6935(
		.A(n_1087),
		.Y(n_1147));

	INVX1 i_6936(
		.A(n_1086),
		.Y(n_1146));

	INVX1 i_6937(
		.A(n_1024),
		.Y(n_931));

	ADDHX1 i_288(
		.A(n_466),
		.B(n_448),
		.S(n_480),
		.CO(n_481));

	ADDHX1 i_289(
		.A(n_467),
		.B(n_449),
		.S(n_482),
		.CO(n_483));

	ADDFHX1 i_290(
		.A(n_431),
		.B(n_413),
		.CI(n_481),
		.S(n_484),
		.CO(n_485));

	ADDHX1 i_291(
		.A(n_468),
		.B(n_450),
		.S(n_486),
		.CO(n_487));

	ADDFHX1 i_292(
		.A(n_432),
		.B(n_414),
		.CI(n_396),
		.S(n_488),
		.CO(n_489));

	ADDFHX1 i_293(
		.A(n_483),
		.B(n_486),
		.CI(n_488),
		.S(n_490),
		.CO(n_491));

	ADDHX1 i_294(
		.A(n_469),
		.B(n_451),
		.S(n_492),
		.CO(n_493));

	ADDFHX1 i_295(
		.A(n_433),
		.B(n_415),
		.CI(n_397),
		.S(n_494),
		.CO(n_495));

	ADDFHX1 i_296(
		.A(n_379),
		.B(n_487),
		.CI(n_489),
		.S(n_496),
		.CO(n_497));

	ADDFHX1 i_297(
		.A(n_492),
		.B(n_494),
		.CI(n_491),
		.S(n_498),
		.CO(n_499));

	ADDHX1 i_298(
		.A(n_470),
		.B(n_452),
		.S(n_500),
		.CO(n_501));

	ADDFHX1 i_299(
		.A(n_434),
		.B(n_416),
		.CI(n_398),
		.S(n_502),
		.CO(n_503));

	ADDFHX1 i_300(
		.A(n_380),
		.B(n_362),
		.CI(n_493),
		.S(n_504),
		.CO(n_505));

	ADDFHX1 i_301(
		.A(n_495),
		.B(n_500),
		.CI(n_502),
		.S(n_506),
		.CO(n_507));

	ADDFHX1 i_302(
		.A(n_497),
		.B(n_504),
		.CI(n_506),
		.S(n_508),
		.CO(n_509));

	ADDHX1 i_303(
		.A(n_471),
		.B(n_453),
		.S(n_510),
		.CO(n_511));

	ADDFHX1 i_304(
		.A(n_435),
		.B(n_417),
		.CI(n_399),
		.S(n_512),
		.CO(n_513));

	ADDFHX1 i_305(
		.A(n_381),
		.B(n_363),
		.CI(n_345),
		.S(n_514),
		.CO(n_515));

	ADDFHX1 i_306(
		.A(n_501),
		.B(n_503),
		.CI(n_510),
		.S(n_516),
		.CO(n_517));

	ADDFHX1 i_307(
		.A(n_512),
		.B(n_514),
		.CI(n_505),
		.S(n_518),
		.CO(n_519));

	ADDFHX1 i_308(
		.A(n_507),
		.B(n_516),
		.CI(n_509),
		.S(n_520),
		.CO(n_521));

	ADDHX1 i_309(
		.A(n_472),
		.B(n_454),
		.S(n_522),
		.CO(n_523));

	ADDFHX1 i_310(
		.A(n_436),
		.B(n_418),
		.CI(n_400),
		.S(n_524),
		.CO(n_525));

	ADDFHX1 i_311(
		.A(n_382),
		.B(n_364),
		.CI(n_346),
		.S(n_526),
		.CO(n_527));

	ADDFHX1 i_312(
		.A(n_328),
		.B(n_511),
		.CI(n_513),
		.S(n_528),
		.CO(n_529));

	ADDFHX1 i_313(
		.A(n_515),
		.B(n_522),
		.CI(n_524),
		.S(n_530),
		.CO(n_531));

	ADDFHX1 i_314(
		.A(n_526),
		.B(n_517),
		.CI(n_528),
		.S(n_532),
		.CO(n_533));

	ADDFHX1 i_315(
		.A(n_530),
		.B(n_519),
		.CI(n_532),
		.S(n_534),
		.CO(n_535));

	ADDHX1 i_316(
		.A(n_473),
		.B(n_455),
		.S(n_536),
		.CO(n_537));

	ADDFHX1 i_317(
		.A(n_437),
		.B(n_419),
		.CI(n_401),
		.S(n_538),
		.CO(n_539));

	ADDFHX1 i_318(
		.A(n_383),
		.B(n_365),
		.CI(n_347),
		.S(n_540),
		.CO(n_541));

	ADDFHX1 i_319(
		.A(n_329),
		.B(n_311),
		.CI(n_523),
		.S(n_542),
		.CO(n_543));

	ADDFHX1 i_320(
		.A(n_525),
		.B(n_527),
		.CI(n_536),
		.S(n_544),
		.CO(n_545));

	ADDFHX1 i_321(
		.A(n_538),
		.B(n_540),
		.CI(n_529),
		.S(n_546),
		.CO(n_547));

	ADDFHX1 i_322(
		.A(n_531),
		.B(n_542),
		.CI(n_544),
		.S(n_548),
		.CO(n_549));

	ADDFHX1 i_323(
		.A(n_533),
		.B(n_546),
		.CI(n_548),
		.S(n_550),
		.CO(n_551));

	ADDHX1 i_324(
		.A(n_474),
		.B(n_456),
		.S(n_552),
		.CO(n_553));

	ADDFHX1 i_325(
		.A(n_438),
		.B(n_420),
		.CI(n_402),
		.S(n_554),
		.CO(n_555));

	ADDFHX1 i_326(
		.A(n_384),
		.B(n_366),
		.CI(n_348),
		.S(n_556),
		.CO(n_557));

	ADDFHX1 i_327(
		.A(n_330),
		.B(n_312),
		.CI(n_294),
		.S(n_558),
		.CO(n_559));

	ADDFHX1 i_328(
		.A(n_537),
		.B(n_539),
		.CI(n_541),
		.S(n_560),
		.CO(n_561));

	ADDFHX1 i_329(
		.A(n_552),
		.B(n_554),
		.CI(n_556),
		.S(n_562),
		.CO(n_563));

	ADDFHX1 i_330(
		.A(n_558),
		.B(n_543),
		.CI(n_545),
		.S(n_564),
		.CO(n_565));

	ADDFHX1 i_331(
		.A(n_560),
		.B(n_562),
		.CI(n_547),
		.S(n_566),
		.CO(n_567));

	ADDFHX1 i_332(
		.A(n_549),
		.B(n_564),
		.CI(n_551),
		.S(n_568),
		.CO(n_569));

	ADDHX1 i_333(
		.A(n_475),
		.B(n_457),
		.S(n_570),
		.CO(n_571));

	ADDFHX1 i_334(
		.A(n_439),
		.B(n_421),
		.CI(n_403),
		.S(n_572),
		.CO(n_573));

	ADDFHX1 i_335(
		.A(n_385),
		.B(n_367),
		.CI(n_349),
		.S(n_574),
		.CO(n_575));

	ADDFHX1 i_336(
		.A(n_331),
		.B(n_313),
		.CI(n_295),
		.S(n_576),
		.CO(n_577));

	ADDFHX1 i_337(
		.A(n_277),
		.B(n_553),
		.CI(n_555),
		.S(n_578),
		.CO(n_579));

	ADDFHX1 i_338(
		.A(n_557),
		.B(n_559),
		.CI(n_570),
		.S(n_580),
		.CO(n_581));

	ADDFHX1 i_339(
		.A(n_572),
		.B(n_574),
		.CI(n_576),
		.S(n_582),
		.CO(n_583));

	ADDFHX1 i_340(
		.A(n_561),
		.B(n_563),
		.CI(n_578),
		.S(n_584),
		.CO(n_585));

	ADDFHX1 i_341(
		.A(n_580),
		.B(n_582),
		.CI(n_565),
		.S(n_586),
		.CO(n_587));

	ADDFHX1 i_342(
		.A(n_584),
		.B(n_567),
		.CI(n_586),
		.S(n_588),
		.CO(n_589));

	ADDHX1 i_343(
		.A(n_476),
		.B(n_458),
		.S(n_590),
		.CO(n_591));

	ADDFHX1 i_344(
		.A(n_440),
		.B(n_422),
		.CI(n_404),
		.S(n_592),
		.CO(n_593));

	ADDFHX1 i_345(
		.A(n_386),
		.B(n_368),
		.CI(n_350),
		.S(n_594),
		.CO(n_595));

	ADDFHX1 i_346(
		.A(n_332),
		.B(n_314),
		.CI(n_296),
		.S(n_596),
		.CO(n_597));

	ADDFHX1 i_347(
		.A(n_278),
		.B(n_260),
		.CI(n_571),
		.S(n_598),
		.CO(n_599));

	ADDFHX1 i_348(
		.A(n_573),
		.B(n_575),
		.CI(n_577),
		.S(n_600),
		.CO(n_601));

	ADDFHX1 i_349(
		.A(n_590),
		.B(n_592),
		.CI(n_594),
		.S(n_602),
		.CO(n_603));

	ADDFHX1 i_350(
		.A(n_596),
		.B(n_579),
		.CI(n_581),
		.S(n_604),
		.CO(n_605));

	ADDFHX1 i_351(
		.A(n_583),
		.B(n_598),
		.CI(n_600),
		.S(n_606),
		.CO(n_607));

	ADDFHX1 i_352(
		.A(n_602),
		.B(n_585),
		.CI(n_604),
		.S(n_608),
		.CO(n_609));

	ADDFHX1 i_353(
		.A(n_606),
		.B(n_587),
		.CI(n_608),
		.S(n_610),
		.CO(n_611));

	ADDHX1 i_354(
		.A(n_477),
		.B(n_459),
		.S(n_612),
		.CO(n_613));

	ADDFHX1 i_355(
		.A(n_441),
		.B(n_423),
		.CI(n_405),
		.S(n_614),
		.CO(n_615));

	ADDFHX1 i_356(
		.A(n_387),
		.B(n_369),
		.CI(n_351),
		.S(n_616),
		.CO(n_617));

	ADDFHX1 i_357(
		.A(n_333),
		.B(n_315),
		.CI(n_297),
		.S(n_618),
		.CO(n_619));

	ADDFHX1 i_358(
		.A(n_279),
		.B(n_261),
		.CI(n_243),
		.S(n_620),
		.CO(n_621));

	ADDFHX1 i_359(
		.A(n_591),
		.B(n_593),
		.CI(n_595),
		.S(n_622),
		.CO(n_623));

	ADDFHX1 i_360(
		.A(n_597),
		.B(n_612),
		.CI(n_614),
		.S(n_624),
		.CO(n_625));

	ADDFHX1 i_361(
		.A(n_616),
		.B(n_618),
		.CI(n_620),
		.S(n_626),
		.CO(n_627));

	ADDFHX1 i_362(
		.A(n_599),
		.B(n_601),
		.CI(n_603),
		.S(n_628),
		.CO(n_629));

	ADDFHX1 i_363(
		.A(n_622),
		.B(n_624),
		.CI(n_626),
		.S(n_630),
		.CO(n_631));

	ADDFHX1 i_364(
		.A(n_605),
		.B(n_607),
		.CI(n_628),
		.S(n_632),
		.CO(n_633));

	ADDFHX1 i_365(
		.A(n_630),
		.B(n_609),
		.CI(n_632),
		.S(n_634),
		.CO(n_635));

	ADDHX1 i_366(
		.A(n_478),
		.B(n_460),
		.S(n_636),
		.CO(n_637));

	ADDFHX1 i_367(
		.A(n_442),
		.B(n_424),
		.CI(n_406),
		.S(n_638),
		.CO(n_639));

	ADDFHX1 i_368(
		.A(n_388),
		.B(n_370),
		.CI(n_352),
		.S(n_640),
		.CO(n_641));

	ADDFHX1 i_369(
		.A(n_334),
		.B(n_316),
		.CI(n_298),
		.S(n_642),
		.CO(n_643));

	ADDFHX1 i_370(
		.A(n_280),
		.B(n_262),
		.CI(n_244),
		.S(n_644),
		.CO(n_645));

	ADDFHX1 i_371(
		.A(n_226),
		.B(n_613),
		.CI(n_615),
		.S(n_646),
		.CO(n_647));

	ADDFHX1 i_372(
		.A(n_617),
		.B(n_619),
		.CI(n_621),
		.S(n_648),
		.CO(n_649));

	ADDFHX1 i_373(
		.A(n_636),
		.B(n_638),
		.CI(n_640),
		.S(n_650),
		.CO(n_651));

	ADDFHX1 i_374(
		.A(n_642),
		.B(n_644),
		.CI(n_623),
		.S(n_652),
		.CO(n_653));

	ADDFHX1 i_375(
		.A(n_625),
		.B(n_627),
		.CI(n_646),
		.S(n_654),
		.CO(n_655));

	ADDFHX1 i_376(
		.A(n_648),
		.B(n_650),
		.CI(n_629),
		.S(n_656),
		.CO(n_657));

	ADDFHX1 i_377(
		.A(n_631),
		.B(n_652),
		.CI(n_654),
		.S(n_658),
		.CO(n_659));

	ADDFHX1 i_378(
		.A(n_633),
		.B(n_656),
		.CI(n_658),
		.S(n_660),
		.CO(n_661));

	ADDHX1 i_379(
		.A(n_479),
		.B(n_461),
		.S(n_662),
		.CO(n_663));

	ADDFHX1 i_380(
		.A(n_443),
		.B(n_425),
		.CI(n_407),
		.S(n_664),
		.CO(n_665));

	ADDFHX1 i_381(
		.A(n_389),
		.B(n_371),
		.CI(n_353),
		.S(n_666),
		.CO(n_667));

	ADDFHX1 i_382(
		.A(n_335),
		.B(n_317),
		.CI(n_299),
		.S(n_668),
		.CO(n_669));

	ADDFHX1 i_383(
		.A(n_281),
		.B(n_263),
		.CI(n_245),
		.S(n_670),
		.CO(n_671));

	ADDFHX1 i_384(
		.A(n_227),
		.B(n_209),
		.CI(n_637),
		.S(n_672),
		.CO(n_673));

	ADDFHX1 i_385(
		.A(n_639),
		.B(n_641),
		.CI(n_643),
		.S(n_674),
		.CO(n_675));

	ADDFHX1 i_386(
		.A(n_645),
		.B(n_662),
		.CI(n_664),
		.S(n_676),
		.CO(n_677));

	ADDFHX1 i_387(
		.A(n_666),
		.B(n_668),
		.CI(n_670),
		.S(n_678),
		.CO(n_679));

	ADDFHX1 i_388(
		.A(n_647),
		.B(n_649),
		.CI(n_651),
		.S(n_680),
		.CO(n_681));

	ADDFHX1 i_389(
		.A(n_672),
		.B(n_674),
		.CI(n_676),
		.S(n_682),
		.CO(n_683));

	ADDFHX1 i_390(
		.A(n_678),
		.B(n_653),
		.CI(n_655),
		.S(n_684),
		.CO(n_685));

	ADDFHX1 i_391(
		.A(n_680),
		.B(n_682),
		.CI(n_657),
		.S(n_686),
		.CO(n_687));

	ADDFHX1 i_392(
		.A(n_659),
		.B(n_684),
		.CI(n_661),
		.S(n_688),
		.CO(n_689));

	ADDHX1 i_393(
		.A(n_462),
		.B(n_444),
		.S(n_690),
		.CO(n_691));

	ADDFHX1 i_394(
		.A(n_426),
		.B(n_408),
		.CI(n_390),
		.S(n_692),
		.CO(n_693));

	ADDFHX1 i_395(
		.A(n_372),
		.B(n_354),
		.CI(n_336),
		.S(n_694),
		.CO(n_695));

	ADDFHX1 i_396(
		.A(n_318),
		.B(n_300),
		.CI(n_282),
		.S(n_696),
		.CO(n_697));

	ADDFHX1 i_397(
		.A(n_264),
		.B(n_246),
		.CI(n_228),
		.S(n_698),
		.CO(n_699));

	ADDFHX1 i_398(
		.A(n_210),
		.B(n_663),
		.CI(n_665),
		.S(n_700),
		.CO(n_701));

	ADDFHX1 i_399(
		.A(n_667),
		.B(n_669),
		.CI(n_671),
		.S(n_702),
		.CO(n_703));

	ADDFHX1 i_400(
		.A(n_690),
		.B(n_692),
		.CI(n_694),
		.S(n_704),
		.CO(n_705));

	ADDFHX1 i_401(
		.A(n_696),
		.B(n_698),
		.CI(n_673),
		.S(n_706),
		.CO(n_707));

	ADDFHX1 i_402(
		.A(n_675),
		.B(n_677),
		.CI(n_679),
		.S(n_708),
		.CO(n_709));

	ADDFHX1 i_403(
		.A(n_700),
		.B(n_702),
		.CI(n_704),
		.S(n_710),
		.CO(n_711));

	ADDFHX1 i_404(
		.A(n_681),
		.B(n_683),
		.CI(n_706),
		.S(n_712),
		.CO(n_713));

	ADDFHX1 i_405(
		.A(n_708),
		.B(n_710),
		.CI(n_685),
		.S(n_714),
		.CO(n_715));

	ADDFHX1 i_406(
		.A(n_712),
		.B(n_687),
		.CI(n_714),
		.S(n_716),
		.CO(n_717));

	ADDFHX1 i_407(
		.A(n_445),
		.B(n_427),
		.CI(n_409),
		.S(n_718),
		.CO(n_719));

	ADDFHX1 i_408(
		.A(n_391),
		.B(n_373),
		.CI(n_355),
		.S(n_720),
		.CO(n_721));

	ADDFHX1 i_409(
		.A(n_337),
		.B(n_319),
		.CI(n_301),
		.S(n_722),
		.CO(n_723));

	ADDFHX1 i_410(
		.A(n_283),
		.B(n_265),
		.CI(n_247),
		.S(n_724),
		.CO(n_725));

	ADDFHX1 i_411(
		.A(n_229),
		.B(n_211),
		.CI(n_691),
		.S(n_726),
		.CO(n_727));

	ADDFHX1 i_412(
		.A(n_693),
		.B(n_695),
		.CI(n_697),
		.S(n_728),
		.CO(n_729));

	ADDFHX1 i_413(
		.A(n_699),
		.B(n_718),
		.CI(n_720),
		.S(n_730),
		.CO(n_731));

	ADDFHX1 i_414(
		.A(n_722),
		.B(n_724),
		.CI(n_701),
		.S(n_732),
		.CO(n_733));

	ADDFHX1 i_415(
		.A(n_703),
		.B(n_705),
		.CI(n_726),
		.S(n_734),
		.CO(n_735));

	ADDFHX1 i_416(
		.A(n_728),
		.B(n_730),
		.CI(n_707),
		.S(n_736),
		.CO(n_737));

	ADDFHX1 i_417(
		.A(n_709),
		.B(n_711),
		.CI(n_732),
		.S(n_738),
		.CO(n_739));

	ADDFHX1 i_418(
		.A(n_734),
		.B(n_713),
		.CI(n_736),
		.S(n_740),
		.CO(n_741));

	ADDFHX1 i_419(
		.A(n_738),
		.B(n_715),
		.CI(n_740),
		.S(n_742),
		.CO(n_743));

	ADDFHX1 i_420(
		.A(n_428),
		.B(n_410),
		.CI(n_392),
		.S(n_744),
		.CO(n_745));

	ADDFHX1 i_421(
		.A(n_374),
		.B(n_356),
		.CI(n_338),
		.S(n_746),
		.CO(n_747));

	ADDFHX1 i_422(
		.A(n_320),
		.B(n_302),
		.CI(n_284),
		.S(n_748),
		.CO(n_749));

	ADDFHX1 i_423(
		.A(n_266),
		.B(n_248),
		.CI(n_230),
		.S(n_750),
		.CO(n_751));

	ADDFHX1 i_424(
		.A(n_212),
		.B(n_719),
		.CI(n_721),
		.S(n_752),
		.CO(n_753));

	ADDFHX1 i_425(
		.A(n_723),
		.B(n_725),
		.CI(n_744),
		.S(n_754),
		.CO(n_755));

	ADDFHX1 i_426(
		.A(n_746),
		.B(n_748),
		.CI(n_750),
		.S(n_756),
		.CO(n_757));

	ADDFHX1 i_427(
		.A(n_727),
		.B(n_729),
		.CI(n_731),
		.S(n_758),
		.CO(n_759));

	ADDFHX1 i_428(
		.A(n_752),
		.B(n_754),
		.CI(n_756),
		.S(n_760),
		.CO(n_761));

	ADDFHX1 i_429(
		.A(n_733),
		.B(n_735),
		.CI(n_758),
		.S(n_762),
		.CO(n_763));

	ADDFHX1 i_430(
		.A(n_760),
		.B(n_737),
		.CI(n_739),
		.S(n_764),
		.CO(n_765));

	ADDFHX1 i_431(
		.A(n_762),
		.B(n_741),
		.CI(n_764),
		.S(n_766),
		.CO(n_767));

	ADDFHX1 i_432(
		.A(n_411),
		.B(n_393),
		.CI(n_375),
		.S(n_768),
		.CO(n_769));

	ADDFHX1 i_433(
		.A(n_357),
		.B(n_339),
		.CI(n_321),
		.S(n_770),
		.CO(n_771));

	ADDFHX1 i_434(
		.A(n_303),
		.B(n_285),
		.CI(n_267),
		.S(n_772),
		.CO(n_773));

	ADDFHX1 i_435(
		.A(n_249),
		.B(n_231),
		.CI(n_213),
		.S(n_774),
		.CO(n_775));

	ADDFHX1 i_436(
		.A(n_745),
		.B(n_747),
		.CI(n_749),
		.S(n_776),
		.CO(n_777));

	ADDFHX1 i_437(
		.A(n_751),
		.B(n_768),
		.CI(n_770),
		.S(n_778),
		.CO(n_779));

	ADDFHX1 i_438(
		.A(n_772),
		.B(n_774),
		.CI(n_753),
		.S(n_780),
		.CO(n_781));

	ADDFHX1 i_439(
		.A(n_755),
		.B(n_757),
		.CI(n_776),
		.S(n_782),
		.CO(n_783));

	ADDFHX1 i_440(
		.A(n_778),
		.B(n_759),
		.CI(n_761),
		.S(n_784),
		.CO(n_785));

	ADDFHX1 i_441(
		.A(n_780),
		.B(n_782),
		.CI(n_763),
		.S(n_786),
		.CO(n_787));

	ADDFHX1 i_442(
		.A(n_784),
		.B(n_765),
		.CI(n_786),
		.S(n_788),
		.CO(n_789));

	ADDFHX1 i_443(
		.A(n_394),
		.B(n_376),
		.CI(n_358),
		.S(n_790),
		.CO(n_791));

	ADDFHX1 i_444(
		.A(n_340),
		.B(n_322),
		.CI(n_304),
		.S(n_792),
		.CO(n_793));

	ADDFHX1 i_445(
		.A(n_286),
		.B(n_268),
		.CI(n_250),
		.S(n_794),
		.CO(n_795));

	ADDFHX1 i_446(
		.A(n_232),
		.B(n_214),
		.CI(n_769),
		.S(n_796),
		.CO(n_797));

	ADDFHX1 i_447(
		.A(n_771),
		.B(n_773),
		.CI(n_775),
		.S(n_798),
		.CO(n_799));

	ADDFHX1 i_448(
		.A(n_790),
		.B(n_792),
		.CI(n_794),
		.S(n_800),
		.CO(n_801));

	ADDFHX1 i_449(
		.A(n_777),
		.B(n_779),
		.CI(n_796),
		.S(n_802),
		.CO(n_803));

	ADDFHX1 i_450(
		.A(n_798),
		.B(n_800),
		.CI(n_781),
		.S(n_804),
		.CO(n_805));

	ADDFHX1 i_451(
		.A(n_783),
		.B(n_802),
		.CI(n_785),
		.S(n_806),
		.CO(n_807));

	ADDFHX1 i_452(
		.A(n_804),
		.B(n_787),
		.CI(n_806),
		.S(n_808),
		.CO(n_809));

	ADDFHX1 i_453(
		.A(n_377),
		.B(n_359),
		.CI(n_341),
		.S(n_810),
		.CO(n_811));

	ADDFHX1 i_454(
		.A(n_323),
		.B(n_305),
		.CI(n_287),
		.S(n_812),
		.CO(n_813));

	ADDFHX1 i_455(
		.A(n_269),
		.B(n_251),
		.CI(n_233),
		.S(n_814),
		.CO(n_815));

	ADDFHX1 i_456(
		.A(n_215),
		.B(n_791),
		.CI(n_793),
		.S(n_816),
		.CO(n_817));

	ADDFHX1 i_457(
		.A(n_795),
		.B(n_810),
		.CI(n_812),
		.S(n_818),
		.CO(n_819));

	ADDFHX1 i_458(
		.A(n_814),
		.B(n_797),
		.CI(n_799),
		.S(n_820),
		.CO(n_821));

	ADDFHX1 i_459(
		.A(n_801),
		.B(n_816),
		.CI(n_818),
		.S(n_822),
		.CO(n_823));

	ADDFHX1 i_460(
		.A(n_803),
		.B(n_820),
		.CI(n_822),
		.S(n_824),
		.CO(n_825));

	ADDFHX1 i_461(
		.A(n_805),
		.B(n_824),
		.CI(n_807),
		.S(n_826),
		.CO(n_827));

	ADDFHX1 i_462(
		.A(n_360),
		.B(n_342),
		.CI(n_324),
		.S(n_828),
		.CO(n_829));

	ADDFHX1 i_463(
		.A(n_306),
		.B(n_288),
		.CI(n_270),
		.S(n_830),
		.CO(n_831));

	ADDFHX1 i_464(
		.A(n_252),
		.B(n_234),
		.CI(n_216),
		.S(n_832),
		.CO(n_833));

	ADDFHX1 i_465(
		.A(n_811),
		.B(n_813),
		.CI(n_815),
		.S(n_834),
		.CO(n_835));

	ADDFHX1 i_466(
		.A(n_828),
		.B(n_830),
		.CI(n_832),
		.S(n_836),
		.CO(n_837));

	ADDFHX1 i_467(
		.A(n_817),
		.B(n_819),
		.CI(n_834),
		.S(n_838),
		.CO(n_839));

	ADDFHX1 i_468(
		.A(n_836),
		.B(n_821),
		.CI(n_823),
		.S(n_840),
		.CO(n_841));

	ADDFHX1 i_469(
		.A(n_838),
		.B(n_825),
		.CI(n_840),
		.S(n_842),
		.CO(n_843));

	ADDFHX1 i_470(
		.A(n_343),
		.B(n_325),
		.CI(n_307),
		.S(n_844),
		.CO(n_845));

	ADDFHX1 i_471(
		.A(n_289),
		.B(n_271),
		.CI(n_253),
		.S(n_846),
		.CO(n_847));

	ADDFHX1 i_472(
		.A(n_235),
		.B(n_217),
		.CI(n_829),
		.S(n_848),
		.CO(n_849));

	ADDFHX1 i_473(
		.A(n_831),
		.B(n_833),
		.CI(n_844),
		.S(n_850),
		.CO(n_851));

	ADDFHX1 i_474(
		.A(n_846),
		.B(n_835),
		.CI(n_837),
		.S(n_852),
		.CO(n_853));

	ADDFHX1 i_475(
		.A(n_848),
		.B(n_850),
		.CI(n_839),
		.S(n_854),
		.CO(n_855));

	ADDFHX1 i_476(
		.A(n_852),
		.B(n_841),
		.CI(n_854),
		.S(n_856),
		.CO(n_857));

	ADDFHX1 i_477(
		.A(n_326),
		.B(n_308),
		.CI(n_290),
		.S(n_858),
		.CO(n_859));

	ADDFHX1 i_478(
		.A(n_272),
		.B(n_254),
		.CI(n_236),
		.S(n_860),
		.CO(n_861));

	ADDFHX1 i_479(
		.A(n_218),
		.B(n_845),
		.CI(n_847),
		.S(n_862),
		.CO(n_863));

	ADDFHX1 i_480(
		.A(n_858),
		.B(n_860),
		.CI(n_849),
		.S(n_864),
		.CO(n_865));

	ADDFHX1 i_481(
		.A(n_851),
		.B(n_862),
		.CI(n_853),
		.S(n_866),
		.CO(n_867));

	ADDFHX1 i_482(
		.A(n_864),
		.B(n_855),
		.CI(n_866),
		.S(n_868),
		.CO(n_869));

	ADDFHX1 i_483(
		.A(n_309),
		.B(n_291),
		.CI(n_273),
		.S(n_870),
		.CO(n_871));

	ADDFHX1 i_484(
		.A(n_255),
		.B(n_237),
		.CI(n_219),
		.S(n_872),
		.CO(n_873));

	ADDFHX1 i_485(
		.A(n_859),
		.B(n_861),
		.CI(n_870),
		.S(n_874),
		.CO(n_875));

	ADDFHX1 i_486(
		.A(n_872),
		.B(n_863),
		.CI(n_874),
		.S(n_876),
		.CO(n_877));

	ADDFHX1 i_487(
		.A(n_865),
		.B(n_876),
		.CI(n_867),
		.S(n_878),
		.CO(n_879));

	ADDFHX1 i_488(
		.A(n_292),
		.B(n_274),
		.CI(n_256),
		.S(n_880),
		.CO(n_881));

	ADDFHX1 i_489(
		.A(n_238),
		.B(n_220),
		.CI(n_871),
		.S(n_882),
		.CO(n_883));

	ADDFHX1 i_490(
		.A(n_873),
		.B(n_880),
		.CI(n_875),
		.S(n_884),
		.CO(n_885));

	ADDFHX1 i_491(
		.A(n_882),
		.B(n_877),
		.CI(n_884),
		.S(n_886),
		.CO(n_887));

	ADDFHX1 i_492(
		.A(n_275),
		.B(n_257),
		.CI(n_239),
		.S(n_888),
		.CO(n_889));

	ADDFHX1 i_493(
		.A(n_221),
		.B(n_881),
		.CI(n_888),
		.S(n_890),
		.CO(n_891));

	ADDFHX1 i_494(
		.A(n_883),
		.B(n_890),
		.CI(n_885),
		.S(n_892),
		.CO(n_893));

	ADDFHX1 i_495(
		.A(n_258),
		.B(n_240),
		.CI(n_222),
		.S(n_894),
		.CO(n_895));

	ADDFHX1 i_496(
		.A(n_889),
		.B(n_894),
		.CI(n_891),
		.S(n_896),
		.CO(n_897));

	ADDFHX1 i_497(
		.A(n_241),
		.B(n_223),
		.CI(n_895),
		.S(n_898),
		.CO(n_899));

	OAI21X1 i_623(
		.A0(n_931),
		.A1(n_901),
		.B0(n_932),
		.Y(n_1025));

	OAI21X1 i_624(
		.A0(n_932),
		.A1(n_902),
		.B0(n_933),
		.Y(n_1026));

	OAI21X1 i_625(
		.A0(n_933),
		.A1(n_903),
		.B0(n_934),
		.Y(n_1027));

	OAI21X1 i_626(
		.A0(n_934),
		.A1(n_904),
		.B0(n_935),
		.Y(n_1028));

	OAI21X1 i_627(
		.A0(n_935),
		.A1(n_905),
		.B0(n_936),
		.Y(n_1029));

	OAI21X1 i_628(
		.A0(n_936),
		.A1(n_906),
		.B0(n_937),
		.Y(n_1030));

	OAI21X1 i_629(
		.A0(n_937),
		.A1(n_907),
		.B0(n_938),
		.Y(n_1031));

	OAI21X1 i_630(
		.A0(n_938),
		.A1(n_908),
		.B0(n_939),
		.Y(n_1032));

	OAI21X1 i_631(
		.A0(n_939),
		.A1(n_909),
		.B0(n_940),
		.Y(n_1033));

	OAI21X1 i_632(
		.A0(n_940),
		.A1(n_910),
		.B0(n_941),
		.Y(n_1034));

	OAI21X1 i_633(
		.A0(n_941),
		.A1(n_911),
		.B0(n_942),
		.Y(n_1035));

	OAI21X1 i_634(
		.A0(n_942),
		.A1(n_912),
		.B0(n_943),
		.Y(n_1036));

	OAI21X1 i_635(
		.A0(n_943),
		.A1(n_913),
		.B0(n_944),
		.Y(n_1037));

	OAI21X1 i_636(
		.A0(n_944),
		.A1(n_914),
		.B0(n_945),
		.Y(n_1038));

	OAI21X1 i_637(
		.A0(n_945),
		.A1(n_915),
		.B0(n_946),
		.Y(n_1039));

	OAI21X1 i_638(
		.A0(n_946),
		.A1(n_916),
		.B0(n_947),
		.Y(n_1040));

	OAI21X1 i_639(
		.A0(n_947),
		.A1(n_917),
		.B0(n_948),
		.Y(n_1041));

	OAI21X1 i_640(
		.A0(n_948),
		.A1(n_918),
		.B0(n_949),
		.Y(n_1042));

	OAI21X1 i_641(
		.A0(n_949),
		.A1(n_919),
		.B0(n_950),
		.Y(n_1043));

	OAI21X1 i_642(
		.A0(n_950),
		.A1(n_920),
		.B0(n_951),
		.Y(n_1044));

	OAI21X1 i_643(
		.A0(n_951),
		.A1(n_921),
		.B0(n_952),
		.Y(n_1045));

	OAI21X1 i_644(
		.A0(n_952),
		.A1(n_922),
		.B0(n_953),
		.Y(n_1046));

	OAI21X1 i_645(
		.A0(n_953),
		.A1(n_923),
		.B0(n_954),
		.Y(n_1047));

	OAI21X1 i_646(
		.A0(n_954),
		.A1(n_924),
		.B0(n_955),
		.Y(n_1048));

	OAI21X1 i_647(
		.A0(n_955),
		.A1(n_925),
		.B0(n_956),
		.Y(n_1049));

	OAI21X1 i_648(
		.A0(n_956),
		.A1(n_926),
		.B0(n_957),
		.Y(n_1050));

	OAI21X1 i_649(
		.A0(n_957),
		.A1(n_927),
		.B0(n_958),
		.Y(n_1051));

	OAI21X1 i_650(
		.A0(n_958),
		.A1(n_928),
		.B0(n_959),
		.Y(n_1052));

	OAI21X1 i_651(
		.A0(n_959),
		.A1(n_929),
		.B0(n_960),
		.Y(n_1053));

	AOI21X1 i_684(
		.A0(n_1024),
		.A1(n_1056),
		.B0(n_1026),
		.Y(n_1086));

	AOI21X1 i_685(
		.A0(n_1025),
		.A1(n_1057),
		.B0(n_1027),
		.Y(n_1087));

	AOI21X1 i_686(
		.A0(n_1026),
		.A1(n_1058),
		.B0(n_1028),
		.Y(n_1088));

	AOI21X1 i_687(
		.A0(n_1027),
		.A1(n_1059),
		.B0(n_1029),
		.Y(n_1089));

	AOI21X1 i_688(
		.A0(n_1028),
		.A1(n_1060),
		.B0(n_1030),
		.Y(n_1090));

	AOI21X1 i_689(
		.A0(n_1029),
		.A1(n_1061),
		.B0(n_1031),
		.Y(n_1091));

	AOI21X1 i_690(
		.A0(n_1030),
		.A1(n_1062),
		.B0(n_1032),
		.Y(n_1092));

	AOI21X1 i_691(
		.A0(n_1031),
		.A1(n_1063),
		.B0(n_1033),
		.Y(n_1093));

	AOI21X1 i_692(
		.A0(n_1032),
		.A1(n_1064),
		.B0(n_1034),
		.Y(n_1094));

	AOI21X1 i_693(
		.A0(n_1033),
		.A1(n_1065),
		.B0(n_1035),
		.Y(n_1095));

	AOI21X1 i_694(
		.A0(n_1034),
		.A1(n_1066),
		.B0(n_1036),
		.Y(n_1096));

	AOI21X1 i_695(
		.A0(n_1035),
		.A1(n_1067),
		.B0(n_1037),
		.Y(n_1097));

	AOI21X1 i_696(
		.A0(n_1036),
		.A1(n_1068),
		.B0(n_1038),
		.Y(n_1098));

	AOI21X1 i_697(
		.A0(n_1037),
		.A1(n_1069),
		.B0(n_1039),
		.Y(n_1099));

	AOI21X1 i_698(
		.A0(n_1038),
		.A1(n_1070),
		.B0(n_1040),
		.Y(n_1100));

	AOI21X1 i_699(
		.A0(n_1039),
		.A1(n_1071),
		.B0(n_1041),
		.Y(n_1101));

	AOI21X1 i_700(
		.A0(n_1040),
		.A1(n_1072),
		.B0(n_1042),
		.Y(n_1102));

	AOI21X1 i_701(
		.A0(n_1041),
		.A1(n_1073),
		.B0(n_1043),
		.Y(n_1103));

	AOI21X1 i_702(
		.A0(n_1042),
		.A1(n_1074),
		.B0(n_1044),
		.Y(n_1104));

	AOI21X1 i_703(
		.A0(n_1043),
		.A1(n_1075),
		.B0(n_1045),
		.Y(n_1105));

	AOI21X1 i_704(
		.A0(n_1044),
		.A1(n_1076),
		.B0(n_1046),
		.Y(n_1106));

	AOI21X1 i_705(
		.A0(n_1045),
		.A1(n_1077),
		.B0(n_1047),
		.Y(n_1107));

	AOI21X1 i_706(
		.A0(n_1046),
		.A1(n_1078),
		.B0(n_1048),
		.Y(n_1108));

	AOI21X1 i_707(
		.A0(n_1047),
		.A1(n_1079),
		.B0(n_1049),
		.Y(n_1109));

	AOI21X1 i_708(
		.A0(n_1048),
		.A1(n_1080),
		.B0(n_1050),
		.Y(n_1110));

	AOI21X1 i_709(
		.A0(n_1049),
		.A1(n_1081),
		.B0(n_1051),
		.Y(n_1111));

	AOI21X1 i_710(
		.A0(n_1050),
		.A1(n_1082),
		.B0(n_1052),
		.Y(n_1112));

	AOI21X1 i_711(
		.A0(n_1051),
		.A1(n_1083),
		.B0(n_1053),
		.Y(n_1113));

	OAI21X1 i_746(
		.A0(n_931),
		.A1(n_1118),
		.B0(n_1088),
		.Y(n_1148));

	OAI21X1 i_747(
		.A0(n_1085),
		.A1(n_1119),
		.B0(n_1089),
		.Y(n_1149));

	OAI21X1 i_748(
		.A0(n_1086),
		.A1(n_1120),
		.B0(n_1090),
		.Y(n_1150));

	OAI21X1 i_749(
		.A0(n_1087),
		.A1(n_1121),
		.B0(n_1091),
		.Y(n_1151));

	OAI21X1 i_750(
		.A0(n_1088),
		.A1(n_1122),
		.B0(n_1092),
		.Y(n_1152));

	OAI21X1 i_751(
		.A0(n_1089),
		.A1(n_1123),
		.B0(n_1093),
		.Y(n_1153));

	OAI21X1 i_752(
		.A0(n_1090),
		.A1(n_1124),
		.B0(n_1094),
		.Y(n_1154));

	OAI21X1 i_753(
		.A0(n_1091),
		.A1(n_1125),
		.B0(n_1095),
		.Y(n_1155));

	OAI21X1 i_754(
		.A0(n_1092),
		.A1(n_1126),
		.B0(n_1096),
		.Y(n_1156));

	OAI21X1 i_755(
		.A0(n_1093),
		.A1(n_1127),
		.B0(n_1097),
		.Y(n_1157));

	OAI21X1 i_756(
		.A0(n_1094),
		.A1(n_1128),
		.B0(n_1098),
		.Y(n_1158));

	OAI21X1 i_757(
		.A0(n_1095),
		.A1(n_1129),
		.B0(n_1099),
		.Y(n_1159));

	OAI21X1 i_758(
		.A0(n_1096),
		.A1(n_1130),
		.B0(n_1100),
		.Y(n_1160));

	OAI21X1 i_759(
		.A0(n_1097),
		.A1(n_1131),
		.B0(n_1101),
		.Y(n_1161));

	OAI21X1 i_760(
		.A0(n_1098),
		.A1(n_1132),
		.B0(n_1102),
		.Y(n_1162));

	OAI21X1 i_761(
		.A0(n_1099),
		.A1(n_1133),
		.B0(n_1103),
		.Y(n_1163));

	OAI21X1 i_762(
		.A0(n_1100),
		.A1(n_1134),
		.B0(n_1104),
		.Y(n_1164));

	OAI21X1 i_763(
		.A0(n_1101),
		.A1(n_1135),
		.B0(n_1105),
		.Y(n_1165));

	OAI21X1 i_764(
		.A0(n_1102),
		.A1(n_1136),
		.B0(n_1106),
		.Y(n_1166));

	OAI21X1 i_765(
		.A0(n_1103),
		.A1(n_1137),
		.B0(n_1107),
		.Y(n_1167));

	OAI21X1 i_766(
		.A0(n_1104),
		.A1(n_1138),
		.B0(n_1108),
		.Y(n_1168));

	OAI21X1 i_767(
		.A0(n_1105),
		.A1(n_1139),
		.B0(n_1109),
		.Y(n_1169));

	OAI21X1 i_768(
		.A0(n_1106),
		.A1(n_1140),
		.B0(n_1110),
		.Y(n_1170));

	OAI21X1 i_769(
		.A0(n_1107),
		.A1(n_1141),
		.B0(n_1111),
		.Y(n_1171));

	OAI21X1 i_770(
		.A0(n_1108),
		.A1(n_1142),
		.B0(n_1112),
		.Y(n_1172));

	OAI21X1 i_771(
		.A0(n_1109),
		.A1(n_1143),
		.B0(n_1113),
		.Y(n_1173));

	AOI21X1 i_810(
		.A0(n_1024),
		.A1(n_1182),
		.B0(n_1152),
		.Y(n_1212));

	AOI21X1 i_811(
		.A0(n_1025),
		.A1(n_1183),
		.B0(n_1153),
		.Y(n_1213));

	AOI21X1 i_812(
		.A0(n_1146),
		.A1(n_1184),
		.B0(n_1154),
		.Y(n_1214));

	AOI21X1 i_813(
		.A0(n_1147),
		.A1(n_1185),
		.B0(n_1155),
		.Y(n_1215));

	AOI21X1 i_814(
		.A0(n_1148),
		.A1(n_1186),
		.B0(n_1156),
		.Y(n_1216));

	AOI21X1 i_815(
		.A0(n_1149),
		.A1(n_1187),
		.B0(n_1157),
		.Y(n_1217));

	AOI21X1 i_816(
		.A0(n_1150),
		.A1(n_1188),
		.B0(n_1158),
		.Y(n_1218));

	AOI21X1 i_817(
		.A0(n_1151),
		.A1(n_1189),
		.B0(n_1159),
		.Y(n_1219));

	AOI21X1 i_818(
		.A0(n_1152),
		.A1(n_1190),
		.B0(n_1160),
		.Y(n_1220));

	AOI21X1 i_819(
		.A0(n_1153),
		.A1(n_1191),
		.B0(n_1161),
		.Y(n_1221));

	AOI21X1 i_820(
		.A0(n_1154),
		.A1(n_1192),
		.B0(n_1162),
		.Y(n_1222));

	AOI21X1 i_821(
		.A0(n_1155),
		.A1(n_1193),
		.B0(n_1163),
		.Y(n_1223));

	AOI21X1 i_822(
		.A0(n_1156),
		.A1(n_1194),
		.B0(n_1164),
		.Y(n_1224));

	AOI21X1 i_823(
		.A0(n_1157),
		.A1(n_1195),
		.B0(n_1165),
		.Y(n_1225));

	AOI21X1 i_824(
		.A0(n_1158),
		.A1(n_1196),
		.B0(n_1166),
		.Y(n_1226));

	AOI21X1 i_825(
		.A0(n_1159),
		.A1(n_1197),
		.B0(n_1167),
		.Y(n_1227));

	AOI21X1 i_826(
		.A0(n_1160),
		.A1(n_1198),
		.B0(n_1168),
		.Y(n_1228));

	AOI21X1 i_827(
		.A0(n_1161),
		.A1(n_1199),
		.B0(n_1169),
		.Y(n_1229));

	AOI21X1 i_828(
		.A0(n_1162),
		.A1(n_1200),
		.B0(n_1170),
		.Y(n_1230));

	AOI21X1 i_829(
		.A0(n_1163),
		.A1(n_1201),
		.B0(n_1171),
		.Y(n_1231));

	AOI21X1 i_830(
		.A0(n_1164),
		.A1(n_1202),
		.B0(n_1172),
		.Y(n_1232));

	AOI21X1 i_831(
		.A0(n_1165),
		.A1(n_1203),
		.B0(n_1173),
		.Y(n_1233));

	OAI21X1 i_878(
		.A0(n_931),
		.A1(n_1250),
		.B0(n_1220),
		.Y(n_1280));

	OAI21X1 i_879(
		.A0(n_1085),
		.A1(n_1251),
		.B0(n_1221),
		.Y(n_1281));

	OAI21X1 i_880(
		.A0(n_1086),
		.A1(n_1252),
		.B0(n_1222),
		.Y(n_1282));

	OAI21X1 i_881(
		.A0(n_1087),
		.A1(n_1253),
		.B0(n_1223),
		.Y(n_1283));

	OAI21X1 i_882(
		.A0(n_1208),
		.A1(n_1254),
		.B0(n_1224),
		.Y(n_1284));

	OAI21X1 i_883(
		.A0(n_1209),
		.A1(n_1255),
		.B0(n_1225),
		.Y(n_1285));

	OAI21X1 i_884(
		.A0(n_1210),
		.A1(n_1256),
		.B0(n_1226),
		.Y(n_1286));

	OAI21X1 i_885(
		.A0(n_1211),
		.A1(n_1257),
		.B0(n_1227),
		.Y(n_1287));

	OAI21X1 i_886(
		.A0(n_1212),
		.A1(n_1258),
		.B0(n_1228),
		.Y(n_1288));

	OAI21X1 i_887(
		.A0(n_1213),
		.A1(n_1259),
		.B0(n_1229),
		.Y(n_1289));

	OAI21X1 i_888(
		.A0(n_1214),
		.A1(n_1260),
		.B0(n_1230),
		.Y(n_1290));

	OAI21X1 i_889(
		.A0(n_1215),
		.A1(n_1261),
		.B0(n_1231),
		.Y(n_1291));

	OAI21X1 i_890(
		.A0(n_1216),
		.A1(n_1262),
		.B0(n_1232),
		.Y(n_1292));

	OAI21X1 i_891(
		.A0(n_1217),
		.A1(n_1263),
		.B0(n_1233),
		.Y(y[31]));

endmodule
module mult_32(
		ovm,
		op_a,
		op_b,
		result);

	input ovm;
	input [15:0] op_a;
	input [15:0] op_b;
	output [31:0] result;




	CLKBUFX3 i_10276(
		.A(n_268),
		.Y(n_7420));

	CLKBUFXL i_10274(
		.A(n_6814),
		.Y(n_7417));

	CLKBUFXL i_10197(
		.A(op_b[0]),
		.Y(n_7307));

	CLKBUFXL i_10187(
		.A(op_a[0]),
		.Y(n_7295));

	BUFX3 i_10163(
		.A(op_b[15]),
		.Y(n_7265));

	BUFX3 i_10160(
		.A(n_7257),
		.Y(n_7260));

	CLKBUFXL i_10157(
		.A(op_a[15]),
		.Y(n_7257));

	CLKBUFXL i_9894(
		.A(n_268),
		.Y(n_6814));

	CLKBUFXL i_9879(
		.A(\ab_a[14] ),
		.Y(n_6789));

	CLKBUFXL i_9878(
		.A(\ab_a[13] ),
		.Y(n_6787));

	CLKBUFXL i_9877(
		.A(\ab_a[12] ),
		.Y(n_6785));

	CLKBUFXL i_9876(
		.A(\ab_a[11] ),
		.Y(n_6783));

	CLKBUFXL i_9875(
		.A(\ab_a[10] ),
		.Y(n_6781));

	CLKBUFXL i_9874(
		.A(\ab_a[9] ),
		.Y(n_6779));

	CLKBUFXL i_9873(
		.A(\ab_a[8] ),
		.Y(n_6777));

	CLKBUFXL i_9872(
		.A(\ab_a[7] ),
		.Y(n_6775));

	CLKBUFXL i_9871(
		.A(\ab_a[6] ),
		.Y(n_6773));

	CLKBUFXL i_9870(
		.A(\ab_a[5] ),
		.Y(n_6771));

	CLKBUFXL i_9869(
		.A(\ab_a[4] ),
		.Y(n_6769));

	CLKBUFXL i_9868(
		.A(\ab_a[3] ),
		.Y(n_6767));

	CLKBUFXL i_9867(
		.A(\ab_a[2] ),
		.Y(n_6765));

	CLKBUFXL i_9866(
		.A(\ab_a[1] ),
		.Y(n_6763));

	CLKBUFXL i_9864(
		.A(\ab_b[14] ),
		.Y(n_6759));

	CLKBUFXL i_9863(
		.A(\ab_b[13] ),
		.Y(n_6757));

	CLKBUFXL i_9862(
		.A(\ab_b[12] ),
		.Y(n_6755));

	CLKBUFXL i_9861(
		.A(\ab_b[11] ),
		.Y(n_6753));

	CLKBUFXL i_9860(
		.A(\ab_b[10] ),
		.Y(n_6751));

	CLKBUFXL i_9859(
		.A(\ab_b[9] ),
		.Y(n_6749));

	CLKBUFXL i_9858(
		.A(\ab_b[8] ),
		.Y(n_6747));

	CLKBUFXL i_9857(
		.A(\ab_b[7] ),
		.Y(n_6745));

	CLKBUFXL i_9856(
		.A(\ab_b[6] ),
		.Y(n_6743));

	CLKBUFXL i_9855(
		.A(\ab_b[5] ),
		.Y(n_6741));

	CLKBUFXL i_9854(
		.A(\ab_b[4] ),
		.Y(n_6739));

	CLKBUFXL i_9853(
		.A(\ab_b[3] ),
		.Y(n_6737));

	CLKBUFXL i_9852(
		.A(\ab_b[2] ),
		.Y(n_6735));

	CLKBUFXL i_9851(
		.A(\ab_b[1] ),
		.Y(n_6733));

	OAI21XL i_818589(
		.A0(\ab_result[22] ),
		.A1(n_588),
		.B0(n_361),
		.Y(result[22]));

	NAND2X1 i_320(
		.A(\ab_result[22] ),
		.B(n_588),
		.Y(n_361));

	OAI21XL i_808588(
		.A0(\ab_result[23] ),
		.A1(n_587),
		.B0(n_359),
		.Y(result[23]));

	NAND2X1 i_317(
		.A(\ab_result[23] ),
		.B(n_587),
		.Y(n_359));

	XOR2X1 i_798587(
		.A(\ab_result[24] ),
		.B(n_586),
		.Y(result[24]));

	OAI21XL i_788586(
		.A0(\ab_result[25] ),
		.A1(n_3099),
		.B0(n_354),
		.Y(result[25]));

	NAND2X1 i_310(
		.A(\ab_result[25] ),
		.B(n_3099),
		.Y(n_354));

	OAI21XL i_778585(
		.A0(\ab_result[26] ),
		.A1(n_584),
		.B0(n_351),
		.Y(result[26]));

	NAND2X1 i_306(
		.A(\ab_result[26] ),
		.B(n_584),
		.Y(n_351));

	OAI21XL i_768584(
		.A0(\ab_result[27] ),
		.A1(n_583),
		.B0(n_348),
		.Y(result[27]));

	NAND2X1 i_302(
		.A(\ab_result[27] ),
		.B(n_583),
		.Y(n_348));

	OAI21XL i_758583(
		.A0(\ab_result[28] ),
		.A1(n_582),
		.B0(n_345),
		.Y(result[28]));

	NAND2X1 i_298(
		.A(\ab_result[28] ),
		.B(n_582),
		.Y(n_345));

	NAND4BXL i_295(
		.AN(n_579),
		.B(n_520),
		.C(n_545),
		.D(n_577),
		.Y(n_344));

	XOR2X1 i_748582(
		.A(\ab_result[29] ),
		.B(n_564),
		.Y(result[29]));

	XOR2X1 i_738581(
		.A(\ab_result[30] ),
		.B(n_549),
		.Y(result[30]));

	OAI21XL i_728580(
		.A0(\ab_result[31] ),
		.A1(n_527),
		.B0(n_336),
		.Y(result[31]));

	NAND2X1 i_250(
		.A(\ab_result[31] ),
		.B(n_527),
		.Y(n_336));

	NOR2BX1 i_238(
		.AN(n_7260),
		.B(n_7265),
		.Y(n_334));

	NOR2BX1 i_237(
		.AN(n_7265),
		.B(n_7260),
		.Y(n_333));

	OAI21XL i_388412(
		.A0(op_b[1]),
		.A1(n_497),
		.B0(n_331),
		.Y(\ab_b[1] ));

	NAND2X1 i_234(
		.A(op_b[1]),
		.B(n_497),
		.Y(n_331));

	OAI21XL i_378411(
		.A0(op_b[2]),
		.A1(n_496),
		.B0(n_329),
		.Y(\ab_b[2] ));

	NAND2X1 i_231(
		.A(op_b[2]),
		.B(n_496),
		.Y(n_329));

	OAI21XL i_368410(
		.A0(op_b[3]),
		.A1(n_495),
		.B0(n_327),
		.Y(\ab_b[3] ));

	NAND2X1 i_228(
		.A(op_b[3]),
		.B(n_495),
		.Y(n_327));

	OAI21XL i_358409(
		.A0(op_b[4]),
		.A1(n_494),
		.B0(n_325),
		.Y(\ab_b[4] ));

	NAND2X1 i_225(
		.A(op_b[4]),
		.B(n_494),
		.Y(n_325));

	OAI21XL i_348408(
		.A0(op_b[5]),
		.A1(n_493),
		.B0(n_322),
		.Y(\ab_b[5] ));

	NAND2X1 i_221(
		.A(op_b[5]),
		.B(n_493),
		.Y(n_322));

	OAI21XL i_338407(
		.A0(op_b[6]),
		.A1(n_492),
		.B0(n_320),
		.Y(\ab_b[6] ));

	NAND2X1 i_218(
		.A(op_b[6]),
		.B(n_492),
		.Y(n_320));

	OAI21XL i_328406(
		.A0(op_b[7]),
		.A1(n_491),
		.B0(n_318),
		.Y(\ab_b[7] ));

	NAND2X1 i_215(
		.A(op_b[7]),
		.B(n_491),
		.Y(n_318));

	OAI21XL i_318405(
		.A0(op_b[8]),
		.A1(n_490),
		.B0(n_316),
		.Y(\ab_b[8] ));

	NAND2X1 i_212(
		.A(op_b[8]),
		.B(n_490),
		.Y(n_316));

	OAI21XL i_308404(
		.A0(op_b[9]),
		.A1(n_489),
		.B0(n_314),
		.Y(\ab_b[9] ));

	NAND2X1 i_209(
		.A(op_b[9]),
		.B(n_489),
		.Y(n_314));

	OAI21XL i_298403(
		.A0(op_b[10]),
		.A1(n_488),
		.B0(n_312),
		.Y(\ab_b[10] ));

	NAND2X1 i_206(
		.A(op_b[10]),
		.B(n_488),
		.Y(n_312));

	OAI21XL i_288402(
		.A0(op_b[11]),
		.A1(n_487),
		.B0(n_310),
		.Y(\ab_b[11] ));

	NAND2X1 i_203(
		.A(op_b[11]),
		.B(n_487),
		.Y(n_310));

	OAI21XL i_278401(
		.A0(op_b[12]),
		.A1(n_486),
		.B0(n_308),
		.Y(\ab_b[12] ));

	NAND2X1 i_200(
		.A(op_b[12]),
		.B(n_486),
		.Y(n_308));

	OAI21XL i_268400(
		.A0(op_b[13]),
		.A1(n_479),
		.B0(n_305),
		.Y(\ab_b[13] ));

	NAND2X1 i_191(
		.A(op_b[13]),
		.B(n_479),
		.Y(n_305));

	OAI21XL i_258399(
		.A0(op_b[14]),
		.A1(n_474),
		.B0(n_302),
		.Y(\ab_b[14] ));

	NAND2X1 i_183(
		.A(op_b[14]),
		.B(n_474),
		.Y(n_302));

	OAI21XL i_388364(
		.A0(op_a[1]),
		.A1(n_451),
		.B0(n_299),
		.Y(\ab_a[1] ));

	NAND2X1 i_168(
		.A(op_a[1]),
		.B(n_451),
		.Y(n_299));

	OAI21XL i_378363(
		.A0(op_a[2]),
		.A1(n_450),
		.B0(n_297),
		.Y(\ab_a[2] ));

	NAND2X1 i_165(
		.A(op_a[2]),
		.B(n_450),
		.Y(n_297));

	OAI21XL i_368362(
		.A0(op_a[3]),
		.A1(n_449),
		.B0(n_295),
		.Y(\ab_a[3] ));

	NAND2X1 i_162(
		.A(op_a[3]),
		.B(n_449),
		.Y(n_295));

	OAI21XL i_358361(
		.A0(op_a[4]),
		.A1(n_448),
		.B0(n_293),
		.Y(\ab_a[4] ));

	NAND2X1 i_159(
		.A(op_a[4]),
		.B(n_448),
		.Y(n_293));

	OAI21XL i_348360(
		.A0(op_a[5]),
		.A1(n_447),
		.B0(n_290),
		.Y(\ab_a[5] ));

	NAND2X1 i_155(
		.A(op_a[5]),
		.B(n_447),
		.Y(n_290));

	OAI21XL i_338359(
		.A0(op_a[6]),
		.A1(n_446),
		.B0(n_288),
		.Y(\ab_a[6] ));

	NAND2X1 i_152(
		.A(op_a[6]),
		.B(n_446),
		.Y(n_288));

	OAI21XL i_328358(
		.A0(op_a[7]),
		.A1(n_445),
		.B0(n_286),
		.Y(\ab_a[7] ));

	NAND2X1 i_142(
		.A(op_a[7]),
		.B(n_445),
		.Y(n_286));

	OAI21XL i_318357(
		.A0(op_a[8]),
		.A1(n_444),
		.B0(n_284),
		.Y(\ab_a[8] ));

	NAND2X1 i_139(
		.A(op_a[8]),
		.B(n_444),
		.Y(n_284));

	OAI21XL i_308356(
		.A0(op_a[9]),
		.A1(n_443),
		.B0(n_282),
		.Y(\ab_a[9] ));

	NAND2X1 i_136(
		.A(op_a[9]),
		.B(n_443),
		.Y(n_282));

	OAI21XL i_298355(
		.A0(op_a[10]),
		.A1(n_442),
		.B0(n_280),
		.Y(\ab_a[10] ));

	NAND2X1 i_133(
		.A(op_a[10]),
		.B(n_442),
		.Y(n_280));

	OAI21XL i_288354(
		.A0(op_a[11]),
		.A1(n_441),
		.B0(n_278),
		.Y(\ab_a[11] ));

	NAND2X1 i_130(
		.A(op_a[11]),
		.B(n_441),
		.Y(n_278));

	OAI21XL i_278353(
		.A0(op_a[12]),
		.A1(n_440),
		.B0(n_276),
		.Y(\ab_a[12] ));

	NAND2X1 i_127(
		.A(op_a[12]),
		.B(n_440),
		.Y(n_276));

	OAI21XL i_268352(
		.A0(op_a[13]),
		.A1(n_433),
		.B0(n_273),
		.Y(\ab_a[13] ));

	NAND2X1 i_118(
		.A(op_a[13]),
		.B(n_433),
		.Y(n_273));

	OAI21XL i_258351(
		.A0(op_a[14]),
		.A1(n_428),
		.B0(n_270),
		.Y(\ab_a[14] ));

	NAND2X1 i_102(
		.A(op_a[14]),
		.B(n_428),
		.Y(n_270));

	NOR2X1 i_6286(
		.A(n_334),
		.B(n_333),
		.Y(n_268));

	OAI21XL i_323(
		.A0(n_558),
		.A1(n_268),
		.B0(\ab_result[21] ),
		.Y(n_363));

	OAI31X1 i_828590(
		.A0(n_7420),
		.A1(\ab_result[21] ),
		.A2(n_558),
		.B0(n_363),
		.Y(result[21]));

	OAI21XL i_326(
		.A0(n_577),
		.A1(n_7417),
		.B0(\ab_result[20] ),
		.Y(n_365));

	OAI31X1 i_838591(
		.A0(n_577),
		.A1(\ab_result[20] ),
		.A2(n_7420),
		.B0(n_365),
		.Y(result[20]));

	OAI21XL i_329(
		.A0(n_515),
		.A1(n_268),
		.B0(\ab_result[19] ),
		.Y(n_367));

	OAI31X1 i_848592(
		.A0(n_7420),
		.A1(\ab_result[19] ),
		.A2(n_515),
		.B0(n_367),
		.Y(result[19]));

	OAI21XL i_332(
		.A0(n_539),
		.A1(n_7417),
		.B0(\ab_result[18] ),
		.Y(n_369));

	OAI31X1 i_858593(
		.A0(n_539),
		.A1(n_7420),
		.A2(\ab_result[18] ),
		.B0(n_369),
		.Y(result[18]));

	XOR2X1 i_868594(
		.A(\ab_result[17] ),
		.B(n_593),
		.Y(result[17]));

	XOR2X1 i_878595(
		.A(\ab_result[16] ),
		.B(n_594),
		.Y(result[16]));

	XOR2X1 i_888596(
		.A(\ab_result[15] ),
		.B(n_595),
		.Y(result[15]));

	XOR2X1 i_898597(
		.A(\ab_result[14] ),
		.B(n_596),
		.Y(result[14]));

	OAI21XL i_347(
		.A0(n_554),
		.A1(n_268),
		.B0(\ab_result[13] ),
		.Y(n_379));

	OAI31X1 i_908598(
		.A0(n_7420),
		.A1(\ab_result[13] ),
		.A2(n_554),
		.B0(n_379),
		.Y(result[13]));

	OAI21XL i_350(
		.A0(n_571),
		.A1(n_7417),
		.B0(\ab_result[12] ),
		.Y(n_381));

	OAI31X1 i_918599(
		.A0(n_571),
		.A1(n_7420),
		.A2(\ab_result[12] ),
		.B0(n_381),
		.Y(result[12]));

	OAI21XL i_353(
		.A0(n_507),
		.A1(n_268),
		.B0(\ab_result[11] ),
		.Y(n_383));

	OAI31X1 i_928600(
		.A0(n_7420),
		.A1(\ab_result[11] ),
		.A2(n_507),
		.B0(n_383),
		.Y(result[11]));

	OAI21XL i_356(
		.A0(n_533),
		.A1(n_268),
		.B0(\ab_result[10] ),
		.Y(n_385));

	OAI31X1 i_938601(
		.A0(n_533),
		.A1(n_7420),
		.A2(\ab_result[10] ),
		.B0(n_385),
		.Y(result[10]));

	NAND2X1 i_359(
		.A(\ab_result[9] ),
		.B(n_601),
		.Y(n_387));

	OAI21XL i_948602(
		.A0(\ab_result[9] ),
		.A1(n_601),
		.B0(n_387),
		.Y(result[9]));

	XOR2X1 i_95(
		.A(\ab_result[8] ),
		.B(n_602),
		.Y(result[8]));

	XOR2X1 i_968603(
		.A(\ab_result[7] ),
		.B(n_603),
		.Y(result[7]));

	XOR2X1 i_97(
		.A(\ab_result[6] ),
		.B(n_604),
		.Y(result[6]));

	XOR2X1 i_98(
		.A(\ab_result[5] ),
		.B(n_605),
		.Y(result[5]));

	NOR2BX1 i_374(
		.AN(n_499),
		.B(\ab_result[3] ),
		.Y(n_397));

	OAI21XL i_375(
		.A0(n_397),
		.A1(n_7417),
		.B0(\ab_result[4] ),
		.Y(n_398));

	OAI31X1 i_998604(
		.A0(n_7420),
		.A1(\ab_result[4] ),
		.A2(n_397),
		.B0(n_398),
		.Y(result[4]));

	OAI21XL i_378(
		.A0(n_499),
		.A1(n_268),
		.B0(\ab_result[3] ),
		.Y(n_400));

	OAI31X1 i_1008605(
		.A0(n_499),
		.A1(n_7420),
		.A2(\ab_result[3] ),
		.B0(n_400),
		.Y(result[3]));

	OAI21XL i_381(
		.A0(n_498),
		.A1(n_7417),
		.B0(\ab_result[2] ),
		.Y(n_402));

	OAI31X1 i_1018606(
		.A0(n_498),
		.A1(n_7420),
		.A2(\ab_result[2] ),
		.B0(n_402),
		.Y(result[2]));

	NAND2X1 i_384(
		.A(\ab_result[1] ),
		.B(n_609),
		.Y(n_404));

	OAI21XL i_1028607(
		.A0(\ab_result[1] ),
		.A1(n_609),
		.B0(n_404),
		.Y(result[1]));

	NOR2X1 i_1(
		.A(op_a[1]),
		.B(op_a[0]),
		.Y(n_406));

	NAND2BX1 i_181705(
		.AN(op_a[2]),
		.B(n_406),
		.Y(n_407));

	NOR2X1 i_39(
		.A(op_a[3]),
		.B(op_a[4]),
		.Y(n_408));

	NOR2X1 i_40(
		.A(op_a[5]),
		.B(op_a[6]),
		.Y(n_409));

	NAND3X1 i_381723(
		.A(n_408),
		.B(n_409),
		.C(n_3101),
		.Y(n_411));

	NOR2X1 i_25(
		.A(op_a[7]),
		.B(op_a[8]),
		.Y(n_412));

	NOR2X1 i_41(
		.A(op_a[9]),
		.B(op_a[10]),
		.Y(n_413));

	NOR4BX1 i_58(
		.AN(n_413),
		.B(op_a[7]),
		.C(op_a[8]),
		.D(n_411),
		.Y(n_415));

	NOR2X1 i_24(
		.A(op_a[11]),
		.B(op_a[12]),
		.Y(n_416));

	NOR2X1 i_89(
		.A(op_a[13]),
		.B(op_a[14]),
		.Y(n_417));

	NOR2X1 i_92(
		.A(op_a[2]),
		.B(op_a[5]),
		.Y(n_420));

	NAND3X1 i_371722(
		.A(n_408),
		.B(n_420),
		.C(n_406),
		.Y(n_422));

	NOR4BX1 i_57(
		.AN(n_412),
		.B(op_a[6]),
		.C(op_a[9]),
		.D(n_422),
		.Y(n_425));

	NOR4X1 i_101(
		.A(op_a[11]),
		.B(op_a[12]),
		.C(op_a[10]),
		.D(op_a[13]),
		.Y(n_427));

	OAI2BB1X1 i_3(
		.A0N(n_425),
		.A1N(n_427),
		.B0(n_7260),
		.Y(n_428));

	NAND2X1 i_361721(
		.A(n_408),
		.B(n_3101),
		.Y(n_429));

	NAND4X1 i_56(
		.A(n_408),
		.B(n_409),
		.C(n_412),
		.D(n_3101),
		.Y(n_431));

	NAND2X1 i_117(
		.A(n_413),
		.B(n_416),
		.Y(n_432));

	OAI21XL i_4(
		.A0(n_431),
		.A1(n_432),
		.B0(n_7260),
		.Y(n_433));

	NOR3X1 i_122(
		.A(op_a[4]),
		.B(op_a[7]),
		.C(op_a[3]),
		.Y(n_435));

	NAND3X1 i_09003(
		.A(n_409),
		.B(n_435),
		.C(n_3101),
		.Y(n_437));

	OR4X1 i_126(
		.A(op_a[9]),
		.B(op_a[10]),
		.C(op_a[8]),
		.D(op_a[11]),
		.Y(n_439));

	OAI21XL i_5(
		.A0(n_437),
		.A1(n_439),
		.B0(n_7257),
		.Y(n_440));

	NAND2BX1 i_42(
		.AN(n_415),
		.B(n_7257),
		.Y(n_441));

	NAND2BX1 i_43(
		.AN(n_425),
		.B(n_7260),
		.Y(n_442));

	NAND2X1 i_44(
		.A(n_7257),
		.B(n_431),
		.Y(n_443));

	NAND2X1 i_45(
		.A(n_7257),
		.B(n_437),
		.Y(n_444));

	NAND2X1 i_46(
		.A(n_7257),
		.B(n_411),
		.Y(n_445));

	NAND2X1 i_47(
		.A(n_7257),
		.B(n_422),
		.Y(n_446));

	NAND2X1 i_48(
		.A(n_7257),
		.B(n_429),
		.Y(n_447));

	OAI21XL i_6(
		.A0(op_a[3]),
		.A1(n_407),
		.B0(op_a[15]),
		.Y(n_448));

	NAND2X1 i_49(
		.A(n_7257),
		.B(n_407),
		.Y(n_449));

	OAI21XL i_50(
		.A0(op_a[1]),
		.A1(op_a[0]),
		.B0(n_7257),
		.Y(n_450));

	NAND2X1 i_51(
		.A(n_7257),
		.B(op_a[0]),
		.Y(n_451));

	NOR2X1 i_11967(
		.A(op_b[1]),
		.B(op_b[0]),
		.Y(n_452));

	NAND2BX1 i_181983(
		.AN(op_b[2]),
		.B(n_452),
		.Y(n_453));

	NOR2X1 i_36(
		.A(op_b[3]),
		.B(op_b[4]),
		.Y(n_454));

	NOR2X1 i_37(
		.A(op_b[5]),
		.B(op_b[6]),
		.Y(n_455));

	NAND3X1 i_382001(
		.A(n_454),
		.B(n_455),
		.C(n_3100),
		.Y(n_457));

	NOR2X1 i_22(
		.A(op_b[7]),
		.B(op_b[8]),
		.Y(n_458));

	NOR2X1 i_38(
		.A(op_b[9]),
		.B(op_b[10]),
		.Y(n_459));

	NOR4BX1 i_582018(
		.AN(n_459),
		.B(op_b[7]),
		.C(op_b[8]),
		.D(n_457),
		.Y(n_461));

	NOR2X1 i_23(
		.A(op_b[11]),
		.B(op_b[12]),
		.Y(n_462));

	NOR2X1 i_173(
		.A(op_b[13]),
		.B(op_b[14]),
		.Y(n_463));

	NOR2X1 i_176(
		.A(op_b[2]),
		.B(op_b[5]),
		.Y(n_466));

	NAND3X1 i_372000(
		.A(n_454),
		.B(n_466),
		.C(n_452),
		.Y(n_468));

	NOR4BX1 i_572017(
		.AN(n_458),
		.B(op_b[6]),
		.C(op_b[9]),
		.D(n_468),
		.Y(n_471));

	NOR4X1 i_182(
		.A(op_b[11]),
		.B(op_b[12]),
		.C(op_b[10]),
		.D(op_b[13]),
		.Y(n_473));

	OAI2BB1X1 i_7(
		.A0N(n_471),
		.A1N(n_473),
		.B0(n_7265),
		.Y(n_474));

	NAND2X1 i_361999(
		.A(n_454),
		.B(n_3100),
		.Y(n_475));

	NAND4X1 i_562016(
		.A(n_454),
		.B(n_455),
		.C(n_458),
		.D(n_3100),
		.Y(n_477));

	NAND2X1 i_190(
		.A(n_459),
		.B(n_462),
		.Y(n_478));

	OAI21XL i_8(
		.A0(n_477),
		.A1(n_478),
		.B0(n_7265),
		.Y(n_479));

	NOR3X1 i_195(
		.A(op_b[4]),
		.B(op_b[7]),
		.C(op_b[3]),
		.Y(n_481));

	NAND3X1 i_2(
		.A(n_455),
		.B(n_481),
		.C(n_3100),
		.Y(n_483));

	OR4X1 i_199(
		.A(op_b[9]),
		.B(op_b[10]),
		.C(op_b[8]),
		.D(op_b[11]),
		.Y(n_485));

	OAI21XL i_9(
		.A0(n_483),
		.A1(n_485),
		.B0(n_7265),
		.Y(n_486));

	NAND2BX1 i_52(
		.AN(n_461),
		.B(n_7265),
		.Y(n_487));

	NAND2BX1 i_53(
		.AN(n_471),
		.B(n_7265),
		.Y(n_488));

	NAND2X1 i_54(
		.A(op_b[15]),
		.B(n_477),
		.Y(n_489));

	NAND2X1 i_55(
		.A(op_b[15]),
		.B(n_483),
		.Y(n_490));

	NAND2X1 i_59(
		.A(n_7265),
		.B(n_457),
		.Y(n_491));

	NAND2X1 i_60(
		.A(op_b[15]),
		.B(n_468),
		.Y(n_492));

	NAND2X1 i_61(
		.A(op_b[15]),
		.B(n_475),
		.Y(n_493));

	OAI21XL i_10(
		.A0(op_b[3]),
		.A1(n_453),
		.B0(op_b[15]),
		.Y(n_494));

	NAND2X1 i_62(
		.A(op_b[15]),
		.B(n_453),
		.Y(n_495));

	OAI21XL i_63(
		.A0(op_b[1]),
		.A1(op_b[0]),
		.B0(op_b[15]),
		.Y(n_496));

	NAND2X1 i_64(
		.A(op_b[15]),
		.B(op_b[0]),
		.Y(n_497));

	NOR2X1 i_12117(
		.A(\ab_result[1] ),
		.B(result[0]),
		.Y(n_498));

	NOR3X1 i_342149(
		.A(\ab_result[1] ),
		.B(result[0]),
		.C(\ab_result[2] ),
		.Y(n_499));

	NOR2X1 i_26(
		.A(\ab_result[3] ),
		.B(\ab_result[4] ),
		.Y(n_500));

	NOR2X1 i_27(
		.A(\ab_result[5] ),
		.B(\ab_result[6] ),
		.Y(n_501));

	NAND3X1 i_702180(
		.A(n_500),
		.B(n_501),
		.C(n_499),
		.Y(n_503));

	NOR2X1 i_28(
		.A(\ab_result[7] ),
		.B(\ab_result[8] ),
		.Y(n_504));

	NOR2X1 i_29(
		.A(\ab_result[9] ),
		.B(\ab_result[10] ),
		.Y(n_505));

	NOR4BX1 i_106(
		.AN(n_505),
		.B(\ab_result[7] ),
		.C(\ab_result[8] ),
		.D(n_503),
		.Y(n_507));

	NOR2X1 i_30(
		.A(\ab_result[11] ),
		.B(\ab_result[12] ),
		.Y(n_508));

	NOR2X1 i_31(
		.A(\ab_result[13] ),
		.B(\ab_result[14] ),
		.Y(n_509));

	NAND3X1 i_110(
		.A(n_508),
		.B(n_509),
		.C(n_507),
		.Y(n_511));

	NOR2X1 i_32(
		.A(\ab_result[15] ),
		.B(\ab_result[16] ),
		.Y(n_512));

	NOR2X1 i_33(
		.A(\ab_result[17] ),
		.B(\ab_result[18] ),
		.Y(n_513));

	NOR4BX1 i_146(
		.AN(n_513),
		.B(\ab_result[15] ),
		.C(\ab_result[16] ),
		.D(n_511),
		.Y(n_515));

	NOR2X1 i_34(
		.A(\ab_result[19] ),
		.B(\ab_result[20] ),
		.Y(n_516));

	NOR2X1 i_35(
		.A(\ab_result[21] ),
		.B(\ab_result[22] ),
		.Y(n_517));

	NAND3X1 i_150(
		.A(n_516),
		.B(n_517),
		.C(n_515),
		.Y(n_519));

	NOR2X1 i_21(
		.A(\ab_result[24] ),
		.B(\ab_result[25] ),
		.Y(n_520));

	OR4X1 i_582170(
		.A(\ab_result[24] ),
		.B(\ab_result[25] ),
		.C(\ab_result[23] ),
		.D(\ab_result[26] ),
		.Y(n_522));

	OR4X1 i_248(
		.A(\ab_result[27] ),
		.B(\ab_result[28] ),
		.C(\ab_result[29] ),
		.D(\ab_result[30] ),
		.Y(n_525));

	OAI32X1 i_11(
		.A0(n_519),
		.A1(n_522),
		.A2(n_525),
		.B0(n_334),
		.B1(n_333),
		.Y(n_527));

	NOR2X1 i_254(
		.A(\ab_result[2] ),
		.B(\ab_result[5] ),
		.Y(n_528));

	NAND3X1 i_692179(
		.A(n_500),
		.B(n_528),
		.C(n_498),
		.Y(n_530));

	NOR4BX1 i_105(
		.AN(n_504),
		.B(\ab_result[6] ),
		.C(\ab_result[9] ),
		.D(n_530),
		.Y(n_533));

	NOR2X1 i_258(
		.A(\ab_result[10] ),
		.B(\ab_result[13] ),
		.Y(n_534));

	NAND3X1 i_109(
		.A(n_508),
		.B(n_534),
		.C(n_533),
		.Y(n_536));

	NOR4BX1 i_145(
		.AN(n_512),
		.B(\ab_result[14] ),
		.C(\ab_result[17] ),
		.D(n_536),
		.Y(n_539));

	NOR4X1 i_263(
		.A(\ab_result[19] ),
		.B(\ab_result[20] ),
		.C(\ab_result[18] ),
		.D(\ab_result[21] ),
		.Y(n_541));

	NAND2X1 i_149(
		.A(n_539),
		.B(n_541),
		.Y(n_542));

	OR4X1 i_572169(
		.A(\ab_result[22] ),
		.B(\ab_result[23] ),
		.C(\ab_result[24] ),
		.D(\ab_result[25] ),
		.Y(n_544));

	NOR2X1 i_20(
		.A(\ab_result[26] ),
		.B(\ab_result[27] ),
		.Y(n_545));

	NOR4BX1 i_267(
		.AN(n_545),
		.B(\ab_result[28] ),
		.C(\ab_result[29] ),
		.D(n_544),
		.Y(n_548));

	AOI31X1 i_12(
		.A0(n_539),
		.A1(n_548),
		.A2(n_541),
		.B0(n_6814),
		.Y(n_549));

	NAND4X1 i_104(
		.A(n_499),
		.B(n_500),
		.C(n_501),
		.D(n_504),
		.Y(n_552));

	NOR4BX1 i_108(
		.AN(n_508),
		.B(\ab_result[9] ),
		.C(\ab_result[10] ),
		.D(n_552),
		.Y(n_554));

	NAND3X1 i_144(
		.A(n_509),
		.B(n_512),
		.C(n_554),
		.Y(n_556));

	NOR4BX1 i_148(
		.AN(n_516),
		.B(\ab_result[17] ),
		.C(\ab_result[18] ),
		.D(n_556),
		.Y(n_558));

	NOR4X1 i_562168(
		.A(\ab_result[21] ),
		.B(\ab_result[22] ),
		.C(\ab_result[23] ),
		.D(\ab_result[24] ),
		.Y(n_560));

	NOR4X1 i_280(
		.A(\ab_result[26] ),
		.B(\ab_result[27] ),
		.C(\ab_result[25] ),
		.D(\ab_result[28] ),
		.Y(n_562));

	AOI31X1 i_13(
		.A0(n_558),
		.A1(n_560),
		.A2(n_562),
		.B0(n_6814),
		.Y(n_564));

	NOR3X1 i_287(
		.A(\ab_result[4] ),
		.B(\ab_result[7] ),
		.C(\ab_result[3] ),
		.Y(n_566));

	NAND3X1 i_712181(
		.A(n_501),
		.B(n_566),
		.C(n_499),
		.Y(n_568));

	NOR4BX1 i_107(
		.AN(n_505),
		.B(\ab_result[8] ),
		.C(\ab_result[11] ),
		.D(n_568),
		.Y(n_571));

	NOR2X1 i_291(
		.A(\ab_result[12] ),
		.B(\ab_result[15] ),
		.Y(n_572));

	NAND3X1 i_111(
		.A(n_509),
		.B(n_572),
		.C(n_571),
		.Y(n_574));

	NOR4BX1 i_147(
		.AN(n_513),
		.B(\ab_result[16] ),
		.C(\ab_result[19] ),
		.D(n_574),
		.Y(n_577));

	NOR2X1 i_285(
		.A(\ab_result[20] ),
		.B(\ab_result[23] ),
		.Y(n_578));

	NAND2X1 i_552167(
		.A(n_517),
		.B(n_578),
		.Y(n_579));

	NAND2BX1 i_14(
		.AN(n_6814),
		.B(n_344),
		.Y(n_582));

	OAI22X1 i_15(
		.A0(n_519),
		.A1(n_522),
		.B0(n_334),
		.B1(n_333),
		.Y(n_583));

	OAI22X1 i_16(
		.A0(n_542),
		.A1(n_544),
		.B0(n_334),
		.B1(n_333),
		.Y(n_584));

	AOI21X1 i_17(
		.A0(n_558),
		.A1(n_560),
		.B0(n_6814),
		.Y(n_585));

	AOI31X1 i_18(
		.A0(n_517),
		.A1(n_578),
		.A2(n_577),
		.B0(n_6814),
		.Y(n_586));

	OAI21XL i_65(
		.A0(n_334),
		.A1(n_333),
		.B0(n_519),
		.Y(n_587));

	OAI21XL i_66(
		.A0(n_334),
		.A1(n_333),
		.B0(n_542),
		.Y(n_588));

	NOR2BX1 i_71(
		.AN(n_556),
		.B(n_6814),
		.Y(n_593));

	NOR2BX1 i_72(
		.AN(n_574),
		.B(n_6814),
		.Y(n_594));

	NOR2BX1 i_73(
		.AN(n_511),
		.B(n_6814),
		.Y(n_595));

	NOR2BX1 i_74(
		.AN(n_536),
		.B(n_6814),
		.Y(n_596));

	OAI21XL i_79(
		.A0(n_334),
		.A1(n_333),
		.B0(n_552),
		.Y(n_601));

	NOR2BX1 i_80(
		.AN(n_568),
		.B(n_6814),
		.Y(n_602));

	NOR2BX1 i_81(
		.AN(n_503),
		.B(n_6814),
		.Y(n_603));

	NOR2BX1 i_82(
		.AN(n_530),
		.B(n_6814),
		.Y(n_604));

	AOI21X1 i_83(
		.A0(n_499),
		.A1(n_500),
		.B0(n_6814),
		.Y(n_605));

	OAI21XL i_86(
		.A0(n_334),
		.A1(n_333),
		.B0(result[0]),
		.Y(n_609));

	AND4X1 i_248350(
		.A(n_416),
		.B(n_417),
		.C(n_7260),
		.D(n_415),
		.Y(\ab_a[15] ));

	AND4X1 i_248398(
		.A(n_462),
		.B(n_463),
		.C(n_7265),
		.D(n_461),
		.Y(\ab_b[15] ));

	INVX1 i_3316(
		.A(n_585),
		.Y(n_3099));

	INVX1 i_3317(
		.A(n_453),
		.Y(n_3100));

	INVX1 i_3318(
		.A(n_407),
		.Y(n_3101));

	m16x16 M16X16_INST(
		.a({
		\ab_a[15] ,
		n_6789,
		n_6787,
		n_6785,
		n_6783,
		n_6781,
		n_6779,
		n_6777,
		n_6775,
		n_6773,
		n_6771,
		n_6769,
		n_6767,
		n_6765,
		n_6763,
		n_7295}),
		.b({
		\ab_b[15] ,
		n_6759,
		n_6757,
		n_6755,
		n_6753,
		n_6751,
		n_6749,
		n_6747,
		n_6745,
		n_6743,
		n_6741,
		n_6739,
		n_6737,
		n_6735,
		n_6733,
		n_7307}),
		.y({
		\ab_result[31] ,
		\ab_result[30] ,
		\ab_result[29] ,
		\ab_result[28] ,
		\ab_result[27] ,
		\ab_result[26] ,
		\ab_result[25] ,
		\ab_result[24] ,
		\ab_result[23] ,
		\ab_result[22] ,
		\ab_result[21] ,
		\ab_result[20] ,
		\ab_result[19] ,
		\ab_result[18] ,
		\ab_result[17] ,
		\ab_result[16] ,
		\ab_result[15] ,
		\ab_result[14] ,
		\ab_result[13] ,
		\ab_result[12] ,
		\ab_result[11] ,
		\ab_result[10] ,
		\ab_result[9] ,
		\ab_result[8] ,
		\ab_result[7] ,
		\ab_result[6] ,
		\ab_result[5] ,
		\ab_result[4] ,
		\ab_result[3] ,
		\ab_result[2] ,
		\ab_result[1] ,
		result[0]}));

endmodule
module port_bus_mach(
		clk,
		reset,
		read,
		write,
		write_h,
		address,
		data_in,
		data_out,
		pad_data_in,
		pad_data_out,
		addrs_in,
		read_cycle,
		sync,
		go,
		as,
		done,
		scan_en,
		BG_scan_in,
		BG_scan_out,
	SPCASCAN_N2_low_mag_8_,
	SPCASCAN_N4_low_mag_3_,
	p_read,
	SPCASCAN_N26_spi_sr_0_,
	FE_PT1_,
	SPCASCAN_N28_read,
	FE_PT2_,
	FE_PT3_,
	SPCASCAN_N29_present_state_1_,
	FE_PT4_,
	FE_PT5_,
	SPCASCAN_N30_ov);
   input SPCASCAN_N2_low_mag_8_;
   input SPCASCAN_N4_low_mag_3_;
   input p_read;
   input SPCASCAN_N26_spi_sr_0_;
   input FE_PT1_;
   output SPCASCAN_N28_read;
   input FE_PT2_;
   input FE_PT3_;
   output SPCASCAN_N29_present_state_1_;
   input FE_PT4_;
   input FE_PT5_;
   input SPCASCAN_N30_ov;

	input clk;
	input reset;
	output read;
	output write;
	output write_h;
	output [2:0] address;
	input [15:0] data_in;
	output [15:0] data_out;
	input [15:0] pad_data_in;
	output [15:0] pad_data_out;
	input [2:0] addrs_in;
	input read_cycle;
	input sync;
	input go;
	output as;
	output done;
	input scan_en;
	input BG_scan_in;
	output BG_scan_out;

	wire [2:0] present_state;



	INVXL i_10648(
		.A(n_7901),
		.Y(BG_scan_out));

	INVXL i_10647(
		.A(write_h),
		.Y(n_7901));

	CLKBUFXL i_10250(
		.A(n_3052),
		.Y(n_7381));

	CLKBUFX3 i_10248(
		.A(n_5006),
		.Y(n_7378));

	INVXL i_9768(
		.A(n_6620),
		.Y(pad_data_out[2]));

	INVXL i_9767(
		.A(data_in[2]),
		.Y(n_6620));

	INVXL i_9765(
		.A(n_6616),
		.Y(pad_data_out[3]));

	INVXL i_9764(
		.A(data_in[3]),
		.Y(n_6616));

	INVXL i_9762(
		.A(n_6612),
		.Y(pad_data_out[4]));

	INVXL i_9761(
		.A(data_in[4]),
		.Y(n_6612));

	INVXL i_9759(
		.A(n_6608),
		.Y(pad_data_out[5]));

	INVXL i_9758(
		.A(data_in[5]),
		.Y(n_6608));

	INVXL i_9756(
		.A(n_6604),
		.Y(pad_data_out[6]));

	INVXL i_9755(
		.A(data_in[6]),
		.Y(n_6604));

	INVXL i_9753(
		.A(n_6600),
		.Y(pad_data_out[7]));

	INVXL i_9752(
		.A(data_in[7]),
		.Y(n_6600));

	INVXL i_9644(
		.A(n_6455),
		.Y(pad_data_out[1]));

	INVXL i_9643(
		.A(data_in[1]),
		.Y(n_6455));

	INVXL i_9623(
		.A(n_6433),
		.Y(pad_data_out[8]));

	INVXL i_9622(
		.A(data_in[8]),
		.Y(n_6433));

	INVXL i_9620(
		.A(n_6429),
		.Y(pad_data_out[9]));

	INVXL i_9619(
		.A(data_in[9]),
		.Y(n_6429));

	INVXL i_9617(
		.A(n_6425),
		.Y(pad_data_out[10]));

	INVXL i_9616(
		.A(data_in[10]),
		.Y(n_6425));

	INVXL i_9614(
		.A(n_6421),
		.Y(pad_data_out[11]));

	INVXL i_9613(
		.A(data_in[11]),
		.Y(n_6421));

	INVXL i_9611(
		.A(n_6417),
		.Y(pad_data_out[12]));

	INVXL i_9610(
		.A(data_in[12]),
		.Y(n_6417));

	INVXL i_9608(
		.A(n_6413),
		.Y(pad_data_out[13]));

	INVXL i_9607(
		.A(data_in[13]),
		.Y(n_6413));

	INVXL i_9605(
		.A(n_6409),
		.Y(pad_data_out[14]));

	INVXL i_9604(
		.A(data_in[14]),
		.Y(n_6409));

	INVXL i_9602(
		.A(n_6405),
		.Y(pad_data_out[15]));

	INVXL i_9601(
		.A(data_in[15]),
		.Y(n_6405));

	CLKBUFXL i_9600(
		.A(addrs_in[0]),
		.Y(address[0]));

	CLKBUFXL i_9597(
		.A(addrs_in[1]),
		.Y(address[1]));

	INVXL i_9593(
		.A(n_6393),
		.Y(address[2]));

	INVXL i_9592(
		.A(addrs_in[2]),
		.Y(n_6393));

	CLKBUFXL i_9504(
		.A(data_in[0]),
		.Y(pad_data_out[0]));

	AOI211X1 i_11(
		.A0(go),
		.A1(read_cycle),
		.B0(SPCASCAN_N29_present_state_1_),
		.C0(present_state[2]),
		.Y(n_11));

	AOI21X1 i_9(
		.A0(present_state[0]),
		.A1(SPCASCAN_N29_present_state_1_),
		.B0(n_3051),
		.Y(n_13));

	NOR4BX1 i_15(
		.AN(go),
		.B(read_cycle),
		.C(present_state[0]),
		.D(SPCASCAN_N29_present_state_1_),
		.Y(n_14));

	OR2X1 i_3(
		.A(n_13),
		.B(n_14),
		.Y(n_15));

	SDFFRHQX1 present_state_reg_0(
		.SI(present_state[2]),
		.SE(scan_en),
		.D(\nbus_616[0] ),
		.CK(clk),
		.RN(n_7381),
		.Q(present_state[0]));

	SDFFRHQX1 present_state_reg_1(
		.SI(BG_scan_out),
		.SE(scan_en),
		.D(n_18),
		.CK(clk),
		.RN(n_7381),
		.Q(SPCASCAN_N29_present_state_1_));

	SDFFRHQX1 present_state_reg_2(
		.SI(done),
		.SE(scan_en),
		.D(n_15),
		.CK(clk),
		.RN(n_7381),
		.Q(present_state[2]));

	SDFFRHQX1 write_reg(
		.SI(present_state[0]),
		.SE(scan_en),
		.D(n_5134),
		.CK(clk),
		.RN(n_7381),
		.Q(write));

	SDFFRHQX1 done_reg(
		.SI(FE_PT2_),
		.SE(scan_en),
		.D(n_5128),
		.CK(clk),
		.RN(n_7381),
		.Q(done));

	SDFFRHQX1 data_out_reg_0(
		.SI(SPCASCAN_N4_low_mag_3_),
		.SE(scan_en),
		.D(n_2949),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[0]));

	MX2X1 i_897(
		.S0(n_7378),
		.B(pad_data_in[0]),
		.A(data_out[0]),
		.Y(n_2949));

	SDFFRHQX1 data_out_reg_1(
		.SI(data_out[2]),
		.SE(scan_en),
		.D(n_2955),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[1]));

	MX2X1 i_904(
		.S0(n_7378),
		.B(pad_data_in[1]),
		.A(data_out[1]),
		.Y(n_2955));

	XOR2X1 i_5(
		.A(SPCASCAN_N29_present_state_1_),
		.B(present_state[0]),
		.Y(n_18));

	SDFFRHQX1 data_out_reg_2(
		.SI(data_out[3]),
		.SE(scan_en),
		.D(n_2961),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[2]));

	MX2X1 i_911(
		.S0(n_7378),
		.B(pad_data_in[2]),
		.A(data_out[2]),
		.Y(n_2961));

	SDFFRHQX1 data_out_reg_3(
		.SI(data_out[6]),
		.SE(scan_en),
		.D(n_2967),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[3]));

	MX2X1 i_918(
		.S0(n_7378),
		.B(pad_data_in[3]),
		.A(data_out[3]),
		.Y(n_2967));

	SDFFRHQX1 data_out_reg_4(
		.SI(SPCASCAN_N2_low_mag_8_),
		.SE(scan_en),
		.D(n_2973),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[4]));

	MX2X1 i_925(
		.S0(n_7378),
		.B(pad_data_in[4]),
		.A(data_out[4]),
		.Y(n_2973));

	OR2X1 i_8(
		.A(n_18),
		.B(n_26),
		.Y(n_21));

	SDFFRHQX1 data_out_reg_5(
		.SI(data_out[4]),
		.SE(scan_en),
		.D(n_2979),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[5]));

	MX2X1 i_932(
		.S0(n_7378),
		.B(pad_data_in[5]),
		.A(data_out[5]),
		.Y(n_2979));

	SDFFRHQX1 data_out_reg_6(
		.SI(p_read),
		.SE(scan_en),
		.D(n_2985),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[6]));

	MX2X1 i_939(
		.S0(n_7378),
		.B(pad_data_in[6]),
		.A(data_out[6]),
		.Y(n_2985));

	SDFFRHQX1 data_out_reg_7(
		.SI(SPCASCAN_N26_spi_sr_0_),
		.SE(scan_en),
		.D(n_2991),
		.CK(clk),
		.RN(n_3052),
		.Q(data_out[7]));

	MX2X1 i_946(
		.S0(n_7378),
		.B(pad_data_in[7]),
		.A(data_out[7]),
		.Y(n_2991));

	SDFFRHQX1 data_out_reg_8(
		.SI(data_out[12]),
		.SE(scan_en),
		.D(n_2997),
		.CK(clk),
		.RN(n_3052),
		.Q(data_out[8]));

	MX2X1 i_953(
		.S0(n_7378),
		.B(pad_data_in[8]),
		.A(data_out[8]),
		.Y(n_2997));

	SDFFRHQX1 data_out_reg_9(
		.SI(FE_PT1_),
		.SE(scan_en),
		.D(n_3003),
		.CK(clk),
		.RN(n_3052),
		.Q(data_out[9]));

	MX2X1 i_960(
		.S0(n_7378),
		.B(pad_data_in[9]),
		.A(data_out[9]),
		.Y(n_3003));

	AOI2BB1X1 i_25(
		.A0N(go),
		.A1N(present_state[2]),
		.B0(SPCASCAN_N29_present_state_1_),
		.Y(n_26));

	SDFFRHQX1 data_out_reg_10(
		.SI(data_out[8]),
		.SE(scan_en),
		.D(n_3009),
		.CK(clk),
		.RN(n_3052),
		.Q(data_out[10]));

	MX2X1 i_967(
		.S0(n_5006),
		.B(pad_data_in[10]),
		.A(data_out[10]),
		.Y(n_3009));

	SDFFRHQX1 data_out_reg_11(
		.SI(data_out[10]),
		.SE(scan_en),
		.D(n_3015),
		.CK(clk),
		.RN(n_3052),
		.Q(data_out[11]));

	MX2X1 i_974(
		.S0(n_7378),
		.B(pad_data_in[11]),
		.A(data_out[11]),
		.Y(n_3015));

	NOR2X1 i_0(
		.A(SPCASCAN_N29_present_state_1_),
		.B(n_3051),
		.Y(n_5134));

	SDFFRHQX1 data_out_reg_12(
		.SI(data_out[9]),
		.SE(scan_en),
		.D(n_3021),
		.CK(clk),
		.RN(n_3052),
		.Q(data_out[12]));

	MX2X1 i_981(
		.S0(n_7378),
		.B(pad_data_in[12]),
		.A(data_out[12]),
		.Y(n_3021));

	AND2X1 i_19001(
		.A(SPCASCAN_N29_present_state_1_),
		.B(present_state[0]),
		.Y(n_5128));

	SDFFRHQX1 data_out_reg_13(
		.SI(FE_PT5_),
		.SE(scan_en),
		.D(n_3027),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[13]));

	MX2X1 i_988(
		.S0(n_7378),
		.B(pad_data_in[13]),
		.A(data_out[13]),
		.Y(n_3027));

	NOR3BX1 i_2(
		.AN(present_state[0]),
		.B(SPCASCAN_N29_present_state_1_),
		.C(present_state[2]),
		.Y(n_5042));

	SDFFRHQX1 data_out_reg_14(
		.SI(data_out[15]),
		.SE(scan_en),
		.D(n_3033),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[14]));

	MX2X1 i_995(
		.S0(n_7378),
		.B(pad_data_in[14]),
		.A(data_out[14]),
		.Y(n_3033));

	NOR2X1 i_7(
		.A(n_11),
		.B(present_state[0]),
		.Y(\nbus_616[0] ));

	SDFFRHQX1 data_out_reg_15(
		.SI(SPCASCAN_N30_ov),
		.SE(scan_en),
		.D(n_3039),
		.CK(clk),
		.RN(n_7381),
		.Q(data_out[15]));

	MX2X1 i_1002(
		.S0(n_7378),
		.B(pad_data_in[15]),
		.A(data_out[15]),
		.Y(n_3039));

	NOR3BX1 i_10(
		.AN(SPCASCAN_N29_present_state_1_),
		.B(present_state[0]),
		.C(present_state[2]),
		.Y(n_5006));

	SDFFRHQX1 read_reg(
		.SI(write),
		.SE(scan_en),
		.D(n_5042),
		.CK(clk),
		.RN(n_3052),
		.Q(SPCASCAN_N28_read));

	SDFFRHQX1 as_reg(
		.SI(FE_PT3_),
		.SE(scan_en),
		.D(n_21),
		.CK(clk),
		.RN(n_3052),
		.Q(as));

	SDFFRHQX1 write_h_reg(
		.SI(FE_PT4_),
		.SE(scan_en),
		.D(n_13),
		.CK(clk),
		.RN(n_3052),
		.Q(write_h));

	INVX1 i_1069(
		.A(present_state[2]),
		.Y(n_3051));

	INVX1 i_1070(
		.A(reset),
		.Y(n_3052));

endmodule
module prog_bus_mach(
		clk,
		reset,
		read,
		write,
		write_h,
		address,
		data_in,
		data_out,
		pad_data_in,
		addrs_in,
		read_cycle,
		sync,
		go,
		as,
		done,
		scan_en,
		BG_scan_in,
		BG_scan_out,
	FE_PT1_,
	FE_PT2_,
	SPCASCAN_N6_present_state_2_,
	FE_PT3_,
	SPCASCAN_N7_present_state_1_,
	FE_PT4_,
	FE_PT5_);
   input FE_PT1_;
   input FE_PT2_;
   output SPCASCAN_N6_present_state_2_;
   input FE_PT3_;
   output SPCASCAN_N7_present_state_1_;
   input FE_PT4_;
   input FE_PT5_;

	input clk;
	input reset;
	output read;
	output write;
	output write_h;
	output [8:0] address;
	input [15:0] data_in;
	output [15:0] data_out;
	input [15:0] pad_data_in;
	input [8:0] addrs_in;
	input read_cycle;
	input sync;
	input go;
	output as;
	output done;
	input scan_en;
	input BG_scan_in;
	output BG_scan_out;

	wire [2:0] present_state;



	INVXL i_10651(
		.A(n_7905),
		.Y(BG_scan_out));

	INVXL i_10650(
		.A(write_h),
		.Y(n_7905));

	CLKBUFXL i_10246(
		.A(n_2937),
		.Y(n_7375));

	CLKBUFX3 i_10244(
		.A(n_4826),
		.Y(n_7372));

	INVXL i_9671(
		.A(n_6491),
		.Y(address[0]));

	INVXL i_9670(
		.A(addrs_in[0]),
		.Y(n_6491));

	INVXL i_9668(
		.A(n_6487),
		.Y(address[1]));

	INVXL i_9667(
		.A(addrs_in[1]),
		.Y(n_6487));

	INVXL i_9665(
		.A(n_6483),
		.Y(address[2]));

	INVXL i_9664(
		.A(addrs_in[2]),
		.Y(n_6483));

	INVXL i_9662(
		.A(n_6479),
		.Y(address[3]));

	INVXL i_9661(
		.A(addrs_in[3]),
		.Y(n_6479));

	INVXL i_9659(
		.A(n_6475),
		.Y(address[4]));

	INVXL i_9658(
		.A(addrs_in[4]),
		.Y(n_6475));

	INVXL i_9656(
		.A(n_6471),
		.Y(address[5]));

	INVXL i_9655(
		.A(addrs_in[5]),
		.Y(n_6471));

	INVXL i_9653(
		.A(n_6467),
		.Y(address[6]));

	INVXL i_9652(
		.A(addrs_in[6]),
		.Y(n_6467));

	INVXL i_9650(
		.A(n_6463),
		.Y(address[7]));

	INVXL i_9649(
		.A(addrs_in[7]),
		.Y(n_6463));

	INVXL i_9647(
		.A(n_6459),
		.Y(address[8]));

	INVXL i_9646(
		.A(addrs_in[8]),
		.Y(n_6459));

	OR3XL i_8(
		.A(n_4835),
		.B(n_20),
		.C(n_18),
		.Y(n_17));

	SDFFRHQX1 present_state_reg_0(
		.SI(as),
		.SE(scan_en),
		.D(\nbus_606[0] ),
		.CK(clk),
		.RN(n_7375),
		.Q(present_state[0]));

	SDFFRHQX1 present_state_reg_1(
		.SI(present_state[0]),
		.SE(scan_en),
		.D(n_20),
		.CK(clk),
		.RN(n_7375),
		.Q(SPCASCAN_N7_present_state_1_));

	SDFFRHQX1 present_state_reg_2(
		.SI(write),
		.SE(scan_en),
		.D(n_21),
		.CK(clk),
		.RN(n_7375),
		.Q(SPCASCAN_N6_present_state_2_));

	SDFFRHQX1 write_reg(
		.SI(done),
		.SE(scan_en),
		.D(n_4954),
		.CK(clk),
		.RN(n_7375),
		.Q(write));

	SDFFRHQX1 data_out_reg_0(
		.SI(data_out[2]),
		.SE(scan_en),
		.D(n_2832),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[0]));

	MX2X1 i_702(
		.S0(n_7372),
		.B(pad_data_in[0]),
		.A(data_out[0]),
		.Y(n_2832));

	NOR2BX1 i_12(
		.AN(go),
		.B(SPCASCAN_N7_present_state_1_),
		.Y(n_18));

	SDFFRHQX1 data_out_reg_1(
		.SI(data_out[15]),
		.SE(scan_en),
		.D(n_2838),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[1]));

	MX2X1 i_709(
		.S0(n_7372),
		.B(pad_data_in[1]),
		.A(data_out[1]),
		.Y(n_2838));

	SDFFRHQX1 data_out_reg_2(
		.SI(data_out[14]),
		.SE(scan_en),
		.D(n_2844),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[2]));

	MX2X1 i_716(
		.S0(n_7372),
		.B(pad_data_in[2]),
		.A(data_out[2]),
		.Y(n_2844));

	XOR2X1 i_5(
		.A(present_state[0]),
		.B(SPCASCAN_N7_present_state_1_),
		.Y(n_20));

	SDFFRHQX1 data_out_reg_3(
		.SI(data_out[4]),
		.SE(scan_en),
		.D(n_2850),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[3]));

	MX2X1 i_723(
		.S0(n_7372),
		.B(pad_data_in[3]),
		.A(data_out[3]),
		.Y(n_2850));

	OAI32X1 i_3(
		.A0(SPCASCAN_N7_present_state_1_),
		.A1(present_state[0]),
		.A2(n_23),
		.B0(n_4868),
		.B1(n_2936),
		.Y(n_21));

	SDFFRHQX1 data_out_reg_4(
		.SI(data_out[8]),
		.SE(scan_en),
		.D(n_2856),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[4]));

	MX2X1 i_730(
		.S0(n_7372),
		.B(pad_data_in[4]),
		.A(data_out[4]),
		.Y(n_2856));

	SDFFRHQX1 data_out_reg_5(
		.SI(data_out[11]),
		.SE(scan_en),
		.D(n_2862),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[5]));

	MX2X1 i_737(
		.S0(n_7372),
		.B(pad_data_in[5]),
		.A(data_out[5]),
		.Y(n_2862));

	NAND2BX1 i_25(
		.AN(read_cycle),
		.B(go),
		.Y(n_23));

	SDFFRHQX1 data_out_reg_6(
		.SI(data_out[0]),
		.SE(scan_en),
		.D(n_2868),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[6]));

	MX2X1 i_744(
		.S0(n_7372),
		.B(pad_data_in[6]),
		.A(data_out[6]),
		.Y(n_2868));

	SDFFRHQX1 data_out_reg_7(
		.SI(data_out[9]),
		.SE(scan_en),
		.D(n_2874),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[7]));

	MX2X1 i_751(
		.S0(n_7372),
		.B(pad_data_in[7]),
		.A(data_out[7]),
		.Y(n_2874));

	AOI21X1 i_21(
		.A0(go),
		.A1(read_cycle),
		.B0(SPCASCAN_N7_present_state_1_),
		.Y(n_25));

	SDFFRHQX1 data_out_reg_8(
		.SI(data_out[7]),
		.SE(scan_en),
		.D(n_2880),
		.CK(clk),
		.RN(n_2937),
		.Q(data_out[8]));

	MX2X1 i_758(
		.S0(n_7372),
		.B(pad_data_in[8]),
		.A(data_out[8]),
		.Y(n_2880));

	SDFFRHQX1 data_out_reg_9(
		.SI(data_out[6]),
		.SE(scan_en),
		.D(n_2886),
		.CK(clk),
		.RN(n_2937),
		.Q(data_out[9]));

	MX2X1 i_765(
		.S0(n_7372),
		.B(pad_data_in[9]),
		.A(data_out[9]),
		.Y(n_2886));

	SDFFRHQX1 data_out_reg_10(
		.SI(data_out[5]),
		.SE(scan_en),
		.D(n_2892),
		.CK(clk),
		.RN(n_2937),
		.Q(data_out[10]));

	MX2X1 i_772(
		.S0(n_4826),
		.B(pad_data_in[10]),
		.A(data_out[10]),
		.Y(n_2892));

	NOR3X1 i_0(
		.A(SPCASCAN_N7_present_state_1_),
		.B(present_state[0]),
		.C(n_2936),
		.Y(n_4954));

	SDFFRHQX1 data_out_reg_11(
		.SI(data_out[12]),
		.SE(scan_en),
		.D(n_2898),
		.CK(clk),
		.RN(n_2937),
		.Q(data_out[11]));

	MX2X1 i_779(
		.S0(n_7372),
		.B(pad_data_in[11]),
		.A(data_out[11]),
		.Y(n_2898));

	AND2X1 i_19000(
		.A(SPCASCAN_N7_present_state_1_),
		.B(present_state[0]),
		.Y(n_4868));

	SDFFRHQX1 data_out_reg_12(
		.SI(FE_PT2_),
		.SE(scan_en),
		.D(n_2904),
		.CK(clk),
		.RN(n_2937),
		.Q(data_out[12]));

	MX2X1 i_786(
		.S0(n_7372),
		.B(pad_data_in[12]),
		.A(data_out[12]),
		.Y(n_2904));

	NOR3BX1 i_2(
		.AN(present_state[0]),
		.B(SPCASCAN_N7_present_state_1_),
		.C(SPCASCAN_N6_present_state_2_),
		.Y(n_4862));

	SDFFRHQX1 data_out_reg_13(
		.SI(FE_PT1_),
		.SE(scan_en),
		.D(n_2910),
		.CK(clk),
		.RN(n_2937),
		.Q(data_out[13]));

	MX2X1 i_793(
		.S0(n_7372),
		.B(pad_data_in[13]),
		.A(data_out[13]),
		.Y(n_2910));

	AOI21X1 i_7(
		.A0(n_25),
		.A1(n_2936),
		.B0(present_state[0]),
		.Y(\nbus_606[0] ));

	SDFFRHQX1 data_out_reg_14(
		.SI(data_out[1]),
		.SE(scan_en),
		.D(n_2916),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[14]));

	MX2X1 i_800(
		.S0(n_7372),
		.B(pad_data_in[14]),
		.A(data_out[14]),
		.Y(n_2916));

	NOR2X1 i_9(
		.A(SPCASCAN_N7_present_state_1_),
		.B(n_2936),
		.Y(n_4835));

	SDFFRHQX1 data_out_reg_15(
		.SI(data_out[10]),
		.SE(scan_en),
		.D(n_2922),
		.CK(clk),
		.RN(n_7375),
		.Q(data_out[15]));

	MX2X1 i_807(
		.S0(n_7372),
		.B(pad_data_in[15]),
		.A(data_out[15]),
		.Y(n_2922));

	NOR3BX1 i_10(
		.AN(SPCASCAN_N7_present_state_1_),
		.B(present_state[0]),
		.C(SPCASCAN_N6_present_state_2_),
		.Y(n_4826));

	SDFFRHQX1 done_reg(
		.SI(FE_PT3_),
		.SE(scan_en),
		.D(n_4868),
		.CK(clk),
		.RN(n_7375),
		.Q(done));

	SDFFRHQX1 read_reg(
		.SI(data_out[3]),
		.SE(scan_en),
		.D(n_4862),
		.CK(clk),
		.RN(n_2937),
		.Q(read));

	SDFFRHQX1 as_reg(
		.SI(FE_PT4_),
		.SE(scan_en),
		.D(n_17),
		.CK(clk),
		.RN(n_2937),
		.Q(as));

	SDFFRHQX1 write_h_reg(
		.SI(FE_PT5_),
		.SE(scan_en),
		.D(n_4835),
		.CK(clk),
		.RN(n_2937),
		.Q(write_h));

	INVX1 i_877(
		.A(SPCASCAN_N6_present_state_2_),
		.Y(n_2936));

	INVX1 i_878(
		.A(reset),
		.Y(n_2937));

endmodule
module tdsp_core_glue(
		addrs_in,
		data_in,
		p_addrs_in,
		p_data_in,
		port_addrs_in,
		port_data_in,
		ar,
		res_adr,
		res_port_adr,
		se_shift_mdr,
		ze_mdr,
		alu_out,
		go_prog,
		read_prog,
		go_data,
		read_data,
		go_port,
		read_port,
		pc_acc,
		arp,
		ar1,
		ar0,
		dp,
		ir,
		pdr,
		opa,
		opb,
		mdr,
		acc,
		pc,
		data_out,
		p_data_out,
		port_data_out,
		top,
		p,
		alu_cmd,
		sel_op_a,
		sel_op_b,
		dec_go_prog,
		enc_go_prog,
		dec_read_prog,
		enc_read_prog,
		dec_go_data,
		enc_go_data,
		dec_read_data,
		enc_read_data,
		dec_go_port,
		enc_go_port,
		dec_read_port,
		enc_read_port,
		dmov_inc);

	output [7:0] addrs_in;
	output [15:0] data_in;
	output [8:0] p_addrs_in;
	output [15:0] p_data_in;
	output [2:0] port_addrs_in;
	output [15:0] port_data_in;
	output [15:0] ar;
	output [7:0] res_adr;
	output [7:0] res_port_adr;
	output [31:0] se_shift_mdr;
	output [31:0] ze_mdr;
	output [15:0] alu_out;
	output go_prog;
	output read_prog;
	output go_data;
	output read_data;
	output go_port;
	output read_port;
	input pc_acc;
	input arp;
	input [15:0] ar1;
	input [15:0] ar0;
	input dp;
	input [15:0] ir;
	output [15:0] pdr;
	output [31:0] opa;
	output [31:0] opb;
	output [15:0] mdr;
	input [32:0] acc;
	input [15:0] pc;
	input [15:0] data_out;
	input [15:0] p_data_out;
	input [15:0] port_data_out;
	input [15:0] top;
	input [31:0] p;
	input [3:0] alu_cmd;
	input [2:0] sel_op_a;
	input [2:0] sel_op_b;
	input dec_go_prog;
	input enc_go_prog;
	input dec_read_prog;
	input enc_read_prog;
	input dec_go_data;
	input enc_go_data;
	input dec_read_data;
	input enc_read_data;
	input dec_go_port;
	input enc_go_port;
	input dec_read_port;
	input enc_read_port;
	input dmov_inc;




	CLKBUFXL i_10414(
		.A(n_1049),
		.Y(n_7604));

	BUFX3 i_10151(
		.A(n_1299),
		.Y(n_7247));

	CLKBUFX3 i_10145(
		.A(n_1359),
		.Y(n_7239));

	BUFX1 i_10142(
		.A(n_1213),
		.Y(n_7236));

	CLKBUFXL i_10139(
		.A(n_402),
		.Y(n_7230));

	BUFX3 i_10137(
		.A(n_410),
		.Y(n_7227));

	BUFXL i_10134(
		.A(n_1357),
		.Y(n_7224));

	CLKBUFXL i_10099(
		.A(n_1041),
		.Y(n_7170));

	BUFX1 i_10097(
		.A(n_1037),
		.Y(n_7167));

	BUFX1 i_10095(
		.A(n_1015),
		.Y(n_7164));

	CLKBUFXL i_10093(
		.A(n_1035),
		.Y(n_7161));

	CLKBUFXL i_10091(
		.A(n_1031),
		.Y(n_7158));

	CLKBUFX3 i_10089(
		.A(n_1023),
		.Y(n_7155));

	CLKBUFX3 i_10087(
		.A(n_1026),
		.Y(n_7152));

	CLKBUFXL i_10055(
		.A(dmov_inc),
		.Y(n_7112));

	CLKBUFXL i_10032(
		.A(n_6255),
		.Y(n_7084));

	CLKBUFX3 i_10021(
		.A(n_1045),
		.Y(n_7060));

	CLKBUFXL i_10019(
		.A(n_1039),
		.Y(n_7056));

	CLKBUFXL i_9997(
		.A(n_1357),
		.Y(n_7015));

	CLKBUFXL i_9992(
		.A(n_1213),
		.Y(n_7006));

	CLKBUFXL i_9990(
		.A(n_1215),
		.Y(n_7003));

	CLKBUFXL i_9989(
		.A(n_1237),
		.Y(n_7001));

	CLKBUFXL i_9967(
		.A(\nbus_686[3] ),
		.Y(opb[3]));

	CLKBUFXL i_9966(
		.A(\nbus_685[2] ),
		.Y(opa[2]));

	CLKBUFXL i_9965(
		.A(\nbus_684[2] ),
		.Y(opb[2]));

	CLKBUFXL i_9963(
		.A(\nbus_683[0] ),
		.Y(opb[0]));

	INVXL i_9833(
		.A(n_6563),
		.Y(mdr[0]));

	INVXL i_9829(
		.A(n_6559),
		.Y(mdr[1]));

	INVXL i_9825(
		.A(n_6555),
		.Y(mdr[2]));

	INVXL i_9821(
		.A(n_6551),
		.Y(mdr[3]));

	INVXL i_9817(
		.A(n_6547),
		.Y(mdr[4]));

	INVXL i_9813(
		.A(n_6543),
		.Y(mdr[5]));

	INVXL i_9809(
		.A(n_6539),
		.Y(mdr[6]));

	INVXL i_9805(
		.A(n_6535),
		.Y(mdr[7]));

	INVXL i_9801(
		.A(n_6531),
		.Y(mdr[8]));

	INVXL i_9797(
		.A(n_6527),
		.Y(mdr[9]));

	INVXL i_9793(
		.A(n_6523),
		.Y(mdr[10]));

	INVXL i_9789(
		.A(n_6519),
		.Y(mdr[11]));

	INVXL i_9785(
		.A(n_6515),
		.Y(mdr[12]));

	INVXL i_9781(
		.A(n_6511),
		.Y(mdr[13]));

	INVXL i_9777(
		.A(n_6507),
		.Y(mdr[14]));

	INVXL i_9773(
		.A(n_6503),
		.Y(mdr[15]));

	INVXL i_9725(
		.A(n_6563),
		.Y(port_data_in[0]));

	INVXL i_9724(
		.A(data_out[0]),
		.Y(n_6563));

	INVXL i_9722(
		.A(n_6559),
		.Y(port_data_in[1]));

	INVXL i_9721(
		.A(data_out[1]),
		.Y(n_6559));

	INVXL i_9719(
		.A(n_6555),
		.Y(port_data_in[2]));

	INVXL i_9718(
		.A(data_out[2]),
		.Y(n_6555));

	INVXL i_9716(
		.A(n_6551),
		.Y(port_data_in[3]));

	INVXL i_9715(
		.A(data_out[3]),
		.Y(n_6551));

	INVXL i_9713(
		.A(n_6547),
		.Y(port_data_in[4]));

	INVXL i_9712(
		.A(data_out[4]),
		.Y(n_6547));

	INVXL i_9710(
		.A(n_6543),
		.Y(port_data_in[5]));

	INVXL i_9709(
		.A(data_out[5]),
		.Y(n_6543));

	INVXL i_9707(
		.A(n_6539),
		.Y(port_data_in[6]));

	INVXL i_9706(
		.A(data_out[6]),
		.Y(n_6539));

	INVXL i_9704(
		.A(n_6535),
		.Y(port_data_in[7]));

	INVXL i_9703(
		.A(data_out[7]),
		.Y(n_6535));

	INVXL i_9701(
		.A(n_6531),
		.Y(port_data_in[8]));

	INVXL i_9700(
		.A(data_out[8]),
		.Y(n_6531));

	INVXL i_9698(
		.A(n_6527),
		.Y(port_data_in[9]));

	INVXL i_9697(
		.A(data_out[9]),
		.Y(n_6527));

	INVXL i_9695(
		.A(n_6523),
		.Y(port_data_in[10]));

	INVXL i_9694(
		.A(data_out[10]),
		.Y(n_6523));

	INVXL i_9692(
		.A(n_6519),
		.Y(port_data_in[11]));

	INVXL i_9691(
		.A(data_out[11]),
		.Y(n_6519));

	INVXL i_9689(
		.A(n_6515),
		.Y(port_data_in[12]));

	INVXL i_9688(
		.A(data_out[12]),
		.Y(n_6515));

	INVXL i_9686(
		.A(n_6511),
		.Y(port_data_in[13]));

	INVXL i_9685(
		.A(data_out[13]),
		.Y(n_6511));

	INVXL i_9683(
		.A(n_6507),
		.Y(port_data_in[14]));

	INVXL i_9682(
		.A(data_out[14]),
		.Y(n_6507));

	INVXL i_9680(
		.A(n_6503),
		.Y(port_data_in[15]));

	INVXL i_9679(
		.A(data_out[15]),
		.Y(n_6503));

	INVX1 i_9677(
		.A(n_6499),
		.Y(port_addrs_in[0]));

	INVXL i_9676(
		.A(ir[8]),
		.Y(n_6499));

	INVX1 i_9674(
		.A(n_6495),
		.Y(port_addrs_in[2]));

	INVXL i_9673(
		.A(ir[10]),
		.Y(n_6495));

	BUFX3 i_9527(
		.A(n_1069),
		.Y(n_6306));

	CLKBUFX3 i_9499(
		.A(arp),
		.Y(n_6255));

	CLKBUFX3 i_9490(
		.A(n_1050),
		.Y(n_6237));

	BUFX3 i_9483(
		.A(ir[9]),
		.Y(port_addrs_in[1]));

	BUFX3 i_9476(
		.A(n_1048),
		.Y(n_6195));

	AOI222X1 i_935(
		.A0(ar0[5]),
		.A1(n_7155),
		.B0(ar1[5]),
		.B1(n_7152),
		.C0(port_data_out[5]),
		.C1(n_7164),
		.Y(n_1100));

	AOI31X1 i_937(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[5]),
		.B0(n_952),
		.Y(n_1097));

	OAI222XL i_939(
		.A0(n_557),
		.A1(n_7604),
		.B0(n_571),
		.B1(n_1086),
		.C0(n_563),
		.C1(n_6237),
		.Y(n_1096));

	AOI22X1 i_941(
		.A0(mdr[4]),
		.A1(n_7112),
		.B0(p_data_out[4]),
		.B1(n_7161),
		.Y(n_1093));

	AOI222X1 i_943(
		.A0(ar0[4]),
		.A1(n_7155),
		.B0(ar1[4]),
		.B1(n_7152),
		.C0(port_data_out[4]),
		.C1(n_7164),
		.Y(n_1092));

	AOI31X1 i_945(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[4]),
		.B0(n_962),
		.Y(n_1089));

	OAI222XL i_947(
		.A0(n_560),
		.A1(n_1049),
		.B0(n_580),
		.B1(n_1086),
		.C0(n_566),
		.C1(n_6237),
		.Y(n_1088));

	NAND3X1 i_33(
		.A(port_addrs_in[2]),
		.B(n_1037),
		.C(port_addrs_in[1]),
		.Y(n_1086));

	AOI22X1 i_949(
		.A0(mdr[3]),
		.A1(n_7112),
		.B0(p_data_out[3]),
		.B1(n_7161),
		.Y(n_1084));

	AOI222X1 i_951(
		.A0(ar0[3]),
		.A1(n_7155),
		.B0(ar1[3]),
		.B1(n_7152),
		.C0(port_data_out[3]),
		.C1(n_7164),
		.Y(n_1083));

	AOI31X1 i_954(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[3]),
		.B0(n_1079),
		.Y(n_1080));

	OAI22X1 i_953(
		.A0(n_571),
		.A1(n_6306),
		.B0(n_570),
		.B1(n_6237),
		.Y(n_1079));

	OAI21XL i_956(
		.A0(n_563),
		.A1(n_7604),
		.B0(n_1077),
		.Y(n_1078));

	AOI22X1 i_955(
		.A0(acc[13]),
		.A1(n_1040),
		.B0(acc[12]),
		.B1(n_1042),
		.Y(n_1077));

	AOI22X1 i_958(
		.A0(mdr[2]),
		.A1(n_7112),
		.B0(p_data_out[2]),
		.B1(n_7161),
		.Y(n_1075));

	AOI222X1 i_960(
		.A0(ar0[2]),
		.A1(n_7155),
		.B0(ar1[2]),
		.B1(n_7152),
		.C0(port_data_out[2]),
		.C1(n_7164),
		.Y(n_1074));

	AOI31X1 i_963(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[2]),
		.B0(n_1070),
		.Y(n_1071));

	OAI22X1 i_962(
		.A0(n_580),
		.A1(n_6306),
		.B0(n_579),
		.B1(n_6237),
		.Y(n_1070));

	OR2X1 i_30(
		.A(port_addrs_in[1]),
		.B(n_1038),
		.Y(n_1069));

	OAI21XL i_965(
		.A0(n_566),
		.A1(n_1049),
		.B0(n_1067),
		.Y(n_1068));

	AOI22X1 i_964(
		.A0(acc[12]),
		.A1(n_1040),
		.B0(acc[11]),
		.B1(n_1042),
		.Y(n_1067));

	AOI22X1 i_967(
		.A0(mdr[1]),
		.A1(n_7112),
		.B0(p_data_out[1]),
		.B1(n_7161),
		.Y(n_1065));

	AOI222X1 i_969(
		.A0(ar0[1]),
		.A1(n_7155),
		.B0(ar1[1]),
		.B1(n_7152),
		.C0(port_data_out[1]),
		.C1(n_7164),
		.Y(n_1064));

	OAI222XL i_972(
		.A0(n_571),
		.A1(n_6237),
		.B0(n_570),
		.B1(n_7604),
		.C0(n_1046),
		.C1(n_4527),
		.Y(n_1061));

	AOI221X1 i_974(
		.A0(acc[10]),
		.A1(n_1042),
		.B0(acc[11]),
		.B1(n_1040),
		.C0(n_997),
		.Y(n_1059));

	AOI22X1 i_976(
		.A0(n_7112),
		.A1(mdr[0]),
		.B0(p_data_out[0]),
		.B1(n_7161),
		.Y(n_1056));

	AOI222X1 i_978(
		.A0(ar0[0]),
		.A1(n_7155),
		.B0(ar1[0]),
		.B1(n_7152),
		.C0(port_data_out[0]),
		.C1(n_7164),
		.Y(n_1055));

	OAI222XL i_981(
		.A0(n_580),
		.A1(n_6237),
		.B0(n_579),
		.B1(n_1049),
		.C0(n_1046),
		.C1(n_4526),
		.Y(n_1052));

	NAND2X1 i_31(
		.A(port_addrs_in[1]),
		.B(n_6195),
		.Y(n_1050));

	NAND2BX1 i_32(
		.AN(port_addrs_in[1]),
		.B(n_6195),
		.Y(n_1049));

	NOR3BX1 i_4(
		.AN(n_1037),
		.B(port_addrs_in[2]),
		.C(n_7060),
		.Y(n_1048));

	NAND2X1 i_9(
		.A(n_7060),
		.B(n_7167),
		.Y(n_1046));

	NOR2X1 i_60(
		.A(n_1013),
		.B(n_1021),
		.Y(n_1045));

	AOI221X1 i_983(
		.A0(acc[9]),
		.A1(n_1042),
		.B0(acc[10]),
		.B1(n_1040),
		.C0(n_1008),
		.Y(n_1044));

	NOR2X1 i_65(
		.A(n_452),
		.B(n_1038),
		.Y(n_1042));

	NOR2X1 i_21(
		.A(ir[8]),
		.B(port_addrs_in[1]),
		.Y(n_1041));

	NOR2X1 i_62(
		.A(n_4506),
		.B(n_1038),
		.Y(n_1040));

	NOR2X1 i_20(
		.A(ir[8]),
		.B(n_4525),
		.Y(n_1039));

	NAND2X1 i_6(
		.A(port_addrs_in[2]),
		.B(n_1037),
		.Y(n_1038));

	NOR4BX1 i_5419(
		.AN(n_1027),
		.B(dmov_inc),
		.C(n_1035),
		.D(n_1015),
		.Y(n_1037));

	NOR4BX1 i_5409(
		.AN(port_addrs_in[2]),
		.B(n_1016),
		.C(n_1030),
		.D(n_1011),
		.Y(n_1035));

	AND2X1 i_22(
		.A(ir[8]),
		.B(n_4525),
		.Y(n_1031));

	NAND3BX1 i_992(
		.AN(ir[12]),
		.B(ir[15]),
		.C(ir[14]),
		.Y(n_1030));

	NOR2X1 i_987(
		.A(n_1026),
		.B(n_1023),
		.Y(n_1027));

	NOR4BBX1 i_5418(
		.AN(n_1020),
		.BN(ir[8]),
		.C(n_1016),
		.D(ir[14]),
		.Y(n_1026));

	NOR4BX1 i_5415(
		.AN(n_1020),
		.B(ir[8]),
		.C(ir[14]),
		.D(n_1016),
		.Y(n_1023));

	NAND2BX1 i_58(
		.AN(ir[8]),
		.B(n_1020),
		.Y(n_1021));

	NOR4BX1 i_16(
		.AN(n_4525),
		.B(port_addrs_in[2]),
		.C(ir[15]),
		.D(n_1017),
		.Y(n_1020));

	NAND2BX1 i_999(
		.AN(ir[11]),
		.B(ir[12]),
		.Y(n_1017));

	NAND2BX1 i_70(
		.AN(dmov_inc),
		.B(ir[13]),
		.Y(n_1016));

	NOR4X1 i_5412(
		.A(ir[15]),
		.B(n_1013),
		.C(ir[12]),
		.D(dmov_inc),
		.Y(n_1015));

	NAND2BX1 i_57(
		.AN(ir[13]),
		.B(ir[14]),
		.Y(n_1013));

	MXI2X1 i_53(
		.S0(ir[11]),
		.B(n_1031),
		.A(n_4508),
		.Y(n_1011));

	NOR2X1 i_666(
		.A(n_578),
		.B(n_1038),
		.Y(n_1008));

	NOR2X1 i_649(
		.A(n_569),
		.B(n_1038),
		.Y(n_997));

	NOR2X1 i_614(
		.A(n_579),
		.B(n_6306),
		.Y(n_962));

	NOR2X1 i_602(
		.A(n_570),
		.B(n_6306),
		.Y(n_952));

	NOR2X1 i_590(
		.A(n_566),
		.B(n_6306),
		.Y(n_942));

	NOR2X1 i_569(
		.A(n_563),
		.B(n_6306),
		.Y(n_932));

	NOR2X1 i_557(
		.A(n_560),
		.B(n_6306),
		.Y(n_922));

	NOR2X1 i_513(
		.A(n_557),
		.B(n_6306),
		.Y(n_912));

	NOR2X1 i_501(
		.A(n_554),
		.B(n_6306),
		.Y(n_902));

	NOR2X1 i_489(
		.A(n_551),
		.B(n_6306),
		.Y(n_892));

	NAND3XL i_453(
		.A(n_1041),
		.B(n_6195),
		.C(acc[30]),
		.Y(n_863));

	NAND3X1 i_442(
		.A(n_7158),
		.B(n_6195),
		.C(acc[30]),
		.Y(n_852));

	NAND3X1 i_441(
		.A(n_1041),
		.B(n_6195),
		.C(acc[31]),
		.Y(n_851));

	NAND3BX1 i_440(
		.AN(n_4506),
		.B(acc[29]),
		.C(n_6195),
		.Y(n_850));

	NOR2BX1 i_581(
		.AN(pc[8]),
		.B(pc_acc),
		.Y(p_addrs_in[8]));

	NAND2X1 i_343(
		.A(mdr[12]),
		.B(n_7003),
		.Y(n_832));

	NAND2X1 i_323(
		.A(p[25]),
		.B(n_7236),
		.Y(n_808));

	NAND2X1 i_13(
		.A(mdr[15]),
		.B(n_1220),
		.Y(n_807));

	NAND2X1 i_315(
		.A(p[24]),
		.B(n_7236),
		.Y(n_799));

	NAND2X1 i_307(
		.A(p[23]),
		.B(n_7236),
		.Y(n_791));

	NAND2X1 i_299(
		.A(p[22]),
		.B(n_7236),
		.Y(n_783));

	NAND2BX1 i_66(
		.AN(n_1221),
		.B(n_1220),
		.Y(n_775));

	AND2X1 i_270(
		.A(n_446),
		.B(n_4507),
		.Y(n_758));

	AND2X1 i_269(
		.A(n_438),
		.B(n_4511),
		.Y(n_757));

	NAND2X1 i_63(
		.A(ir[12]),
		.B(n_4504),
		.Y(n_719));

	NOR2X1 i_208(
		.A(n_1314),
		.B(n_1218),
		.Y(n_701));

	NAND2X1 i_181(
		.A(ir[7]),
		.B(n_4504),
		.Y(n_672));

	NAND2X1 i_176(
		.A(ir[6]),
		.B(n_4504),
		.Y(n_667));

	NAND2X1 i_169(
		.A(n_1308),
		.B(n_4507),
		.Y(n_660));

	NAND2X1 i_166(
		.A(ir[4]),
		.B(n_4504),
		.Y(n_657));

	NAND2X1 i_89(
		.A(top[3]),
		.B(n_7239),
		.Y(n_604));

	NAND2X1 i_85(
		.A(top[2]),
		.B(n_7239),
		.Y(n_600));

	NAND2X1 i_77(
		.A(top[0]),
		.B(n_7239),
		.Y(n_592));

	MXI2X1 i_152250(
		.S0(port_addrs_in[0]),
		.B(acc[13]),
		.A(acc[14]),
		.Y(n_580));

	MXI2X1 i_172252(
		.S0(port_addrs_in[0]),
		.B(acc[15]),
		.A(acc[16]),
		.Y(n_579));

	AOI22X1 i_72(
		.A0(acc[12]),
		.A1(n_1041),
		.B0(acc[11]),
		.B1(n_1031),
		.Y(n_578));

	MXI2X1 i_162251(
		.S0(port_addrs_in[0]),
		.B(acc[14]),
		.A(acc[15]),
		.Y(n_571));

	MXI2X1 i_182253(
		.S0(port_addrs_in[0]),
		.B(acc[16]),
		.A(acc[17]),
		.Y(n_570));

	AOI22X1 i_73(
		.A0(acc[13]),
		.A1(n_1041),
		.B0(acc[12]),
		.B1(n_1031),
		.Y(n_569));

	MXI2X1 i_192254(
		.S0(port_addrs_in[0]),
		.B(acc[17]),
		.A(acc[18]),
		.Y(n_566));

	MXI2X1 i_202255(
		.S0(port_addrs_in[0]),
		.B(acc[18]),
		.A(acc[19]),
		.Y(n_563));

	MXI2X1 i_212256(
		.S0(port_addrs_in[0]),
		.B(acc[19]),
		.A(acc[20]),
		.Y(n_560));

	MXI2X1 i_222257(
		.S0(port_addrs_in[0]),
		.B(acc[20]),
		.A(acc[21]),
		.Y(n_557));

	MXI2X1 i_23(
		.S0(port_addrs_in[0]),
		.B(acc[21]),
		.A(acc[22]),
		.Y(n_554));

	MXI2X1 i_242258(
		.S0(port_addrs_in[0]),
		.B(acc[22]),
		.A(acc[23]),
		.Y(n_551));

	MXI2X1 i_252259(
		.S0(ir[8]),
		.B(acc[23]),
		.A(acc[24]),
		.Y(n_548));

	MXI2X1 i_262260(
		.S0(ir[8]),
		.B(acc[24]),
		.A(acc[25]),
		.Y(n_545));

	MXI2X1 i_272261(
		.S0(port_addrs_in[0]),
		.B(acc[25]),
		.A(acc[26]),
		.Y(n_542));

	MXI2X1 i_282262(
		.S0(port_addrs_in[0]),
		.B(acc[26]),
		.A(acc[27]),
		.Y(n_539));

	NAND2X1 i_390(
		.A(n_1208),
		.B(n_1194),
		.Y(n_489));

	NAND2X1 i_388(
		.A(n_1207),
		.B(n_1195),
		.Y(n_487));

	NAND2X1 i_386(
		.A(n_1206),
		.B(n_1196),
		.Y(n_485));

	NAND2X1 i_384(
		.A(n_1205),
		.B(n_1197),
		.Y(n_483));

	NAND2X1 i_383(
		.A(n_1204),
		.B(n_1198),
		.Y(n_482));

	NAND2X1 i_381(
		.A(n_1210),
		.B(n_1199),
		.Y(n_480));

	NAND2X1 i_379(
		.A(n_1209),
		.B(n_1201),
		.Y(n_478));

	AOI21X1 i_74(
		.A0(sel_op_b[0]),
		.A1(sel_op_b[1]),
		.B0(sel_op_b[2]),
		.Y(n_456));

	NAND2X1 i_75(
		.A(ir[8]),
		.B(port_addrs_in[1]),
		.Y(n_452));

	AOI22X1 i_51(
		.A0(mdr[14]),
		.A1(n_4508),
		.B0(mdr[15]),
		.B1(n_452),
		.Y(n_449));

	AOI222X1 i_50(
		.A0(mdr[13]),
		.A1(n_4508),
		.B0(mdr[14]),
		.B1(n_7056),
		.C0(mdr[15]),
		.C1(n_4525),
		.Y(n_447));

	NAND2X1 i_49(
		.A(n_1228),
		.B(n_1227),
		.Y(n_446));

	NAND2X1 i_48(
		.A(n_1232),
		.B(n_1231),
		.Y(n_445));

	NAND2X1 i_47(
		.A(n_1236),
		.B(n_1235),
		.Y(n_444));

	AOI221XL i_46(
		.A0(mdr[9]),
		.A1(n_4508),
		.B0(mdr[10]),
		.B1(n_7056),
		.C0(n_4510),
		.Y(n_443));

	NAND2X1 i_45(
		.A(n_1247),
		.B(n_1246),
		.Y(n_442));

	NAND2X1 i_44(
		.A(n_1252),
		.B(n_1251),
		.Y(n_441));

	NAND2X1 i_43(
		.A(n_1257),
		.B(n_1256),
		.Y(n_440));

	NAND2X1 i_42(
		.A(n_1264),
		.B(n_1263),
		.Y(n_439));

	NAND2X1 i_41(
		.A(n_1270),
		.B(n_1269),
		.Y(n_438));

	NAND2X1 i_40(
		.A(n_1276),
		.B(n_1275),
		.Y(n_437));

	NAND2X1 i_39(
		.A(n_1282),
		.B(n_1281),
		.Y(n_436));

	NAND2X1 i_38(
		.A(n_1289),
		.B(n_1288),
		.Y(n_435));

	MXI2X1 i_22222(
		.S0(port_addrs_in[0]),
		.B(mdr[0]),
		.A(mdr[1]),
		.Y(n_432));

	OAI21XL i_37(
		.A0(n_432),
		.A1(n_4525),
		.B0(n_1294),
		.Y(n_430));

	AOI222X1 i_36(
		.A0(mdr[2]),
		.A1(n_1041),
		.B0(mdr[1]),
		.B1(n_7158),
		.C0(mdr[0]),
		.C1(n_7056),
		.Y(n_428));

	OAI21XL i_09007(
		.A0(sel_op_a[1]),
		.A1(n_4520),
		.B0(sel_op_a[0]),
		.Y(n_410));

	NAND2X1 i_7(
		.A(mdr[15]),
		.B(n_7227),
		.Y(n_402));

	AOI22X1 i_933(
		.A0(mdr[5]),
		.A1(n_7112),
		.B0(p_data_out[5]),
		.B1(n_7161),
		.Y(n_1101));

	OAI222XL i_931(
		.A0(n_554),
		.A1(n_7604),
		.B0(n_579),
		.B1(n_1086),
		.C0(n_560),
		.C1(n_6237),
		.Y(n_1104));

	AOI31X1 i_929(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[6]),
		.B0(n_942),
		.Y(n_1105));

	AOI222X1 i_927(
		.A0(ar0[6]),
		.A1(n_7155),
		.B0(ar1[6]),
		.B1(n_7152),
		.C0(port_data_out[6]),
		.C1(n_7164),
		.Y(n_1108));

	AOI22X1 i_925(
		.A0(mdr[6]),
		.A1(n_7112),
		.B0(p_data_out[6]),
		.B1(n_7161),
		.Y(n_1109));

	OAI222XL i_923(
		.A0(n_551),
		.A1(n_7604),
		.B0(n_570),
		.B1(n_1086),
		.C0(n_557),
		.C1(n_6237),
		.Y(n_1112));

	AOI31X1 i_921(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[7]),
		.B0(n_932),
		.Y(n_1113));

	AOI222X1 i_919(
		.A0(ar0[7]),
		.A1(n_7155),
		.B0(ar1[7]),
		.B1(n_7152),
		.C0(port_data_out[7]),
		.C1(n_7164),
		.Y(n_1116));

	AOI22X1 i_917(
		.A0(mdr[7]),
		.A1(n_7112),
		.B0(p_data_out[7]),
		.B1(n_7161),
		.Y(n_1117));

	OAI222XL i_915(
		.A0(n_548),
		.A1(n_1049),
		.B0(n_566),
		.B1(n_1086),
		.C0(n_554),
		.C1(n_6237),
		.Y(n_1120));

	AOI31X1 i_913(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[8]),
		.B0(n_922),
		.Y(n_1121));

	AOI222X1 i_911(
		.A0(ar0[8]),
		.A1(n_7155),
		.B0(ar1[8]),
		.B1(n_7152),
		.C0(port_data_out[8]),
		.C1(n_7164),
		.Y(n_1124));

	AOI22X1 i_909(
		.A0(mdr[8]),
		.A1(n_7112),
		.B0(p_data_out[8]),
		.B1(n_7161),
		.Y(n_1125));

	OAI222XL i_907(
		.A0(n_545),
		.A1(n_7604),
		.B0(n_563),
		.B1(n_1086),
		.C0(n_551),
		.C1(n_6237),
		.Y(n_1128));

	AOI31X1 i_905(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[9]),
		.B0(n_912),
		.Y(n_1129));

	AOI222X1 i_903(
		.A0(ar0[9]),
		.A1(n_7155),
		.B0(ar1[9]),
		.B1(n_7152),
		.C0(port_data_out[9]),
		.C1(n_7164),
		.Y(n_1132));

	AOI22X1 i_901(
		.A0(mdr[9]),
		.A1(n_7112),
		.B0(p_data_out[9]),
		.B1(n_7161),
		.Y(n_1133));

	OAI222XL i_899(
		.A0(n_542),
		.A1(n_1049),
		.B0(n_560),
		.B1(n_1086),
		.C0(n_548),
		.C1(n_6237),
		.Y(n_1136));

	AOI31X1 i_897(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[10]),
		.B0(n_902),
		.Y(n_1137));

	AOI222X1 i_895(
		.A0(ar0[10]),
		.A1(n_7155),
		.B0(ar1[10]),
		.B1(n_7152),
		.C0(port_data_out[10]),
		.C1(n_7164),
		.Y(n_1140));

	AOI22X1 i_893(
		.A0(mdr[10]),
		.A1(n_7112),
		.B0(p_data_out[10]),
		.B1(n_7161),
		.Y(n_1141));

	OAI222XL i_891(
		.A0(n_539),
		.A1(n_1049),
		.B0(n_557),
		.B1(n_1086),
		.C0(n_545),
		.C1(n_6237),
		.Y(n_1144));

	AOI31X1 i_889(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[11]),
		.B0(n_892),
		.Y(n_1145));

	AOI222X1 i_887(
		.A0(ar0[11]),
		.A1(n_7155),
		.B0(ar1[11]),
		.B1(n_7152),
		.C0(port_data_out[11]),
		.C1(n_7164),
		.Y(n_1148));

	AOI22X1 i_885(
		.A0(mdr[11]),
		.A1(n_7112),
		.B0(p_data_out[11]),
		.B1(n_7161),
		.Y(n_1149));

	NAND2X1 i_61(
		.A(acc[28]),
		.B(n_6195),
		.Y(n_1152));

	AOI32X1 i_882(
		.A0(n_1031),
		.A1(n_6195),
		.A2(acc[27]),
		.B0(n_1041),
		.B1(n_4514),
		.Y(n_1153));

	OAI21XL i_883(
		.A0(n_554),
		.A1(n_1086),
		.B0(n_1153),
		.Y(n_1154));

	OAI22X1 i_880(
		.A0(n_548),
		.A1(n_6306),
		.B0(n_542),
		.B1(n_6237),
		.Y(n_1155));

	AOI31X1 i_881(
		.A0(n_7060),
		.A1(n_7167),
		.A2(acc[12]),
		.B0(n_1155),
		.Y(n_1156));

	AOI222X1 i_878(
		.A0(ar0[12]),
		.A1(n_7155),
		.B0(ar1[12]),
		.B1(n_7152),
		.C0(port_data_out[12]),
		.C1(n_7164),
		.Y(n_1159));

	AOI22X1 i_876(
		.A0(mdr[12]),
		.A1(n_7112),
		.B0(p_data_out[12]),
		.B1(n_7161),
		.Y(n_1160));

	AOI32X1 i_873(
		.A0(n_1041),
		.A1(n_6195),
		.A2(acc[29]),
		.B0(n_1031),
		.B1(n_4514),
		.Y(n_1163));

	OAI21XL i_874(
		.A0(n_551),
		.A1(n_1086),
		.B0(n_1163),
		.Y(n_1164));

	OAI22X1 i_871(
		.A0(n_545),
		.A1(n_6306),
		.B0(n_539),
		.B1(n_6237),
		.Y(n_1165));

	AOI31X1 i_872(
		.A0(n_7060),
		.A1(acc[13]),
		.A2(n_7167),
		.B0(n_1165),
		.Y(n_1166));

	AOI222X1 i_869(
		.A0(ar0[13]),
		.A1(n_7155),
		.B0(ar1[13]),
		.B1(n_7152),
		.C0(port_data_out[13]),
		.C1(n_7164),
		.Y(n_1169));

	AOI22X1 i_867(
		.A0(mdr[13]),
		.A1(n_7112),
		.B0(p_data_out[13]),
		.B1(n_7161),
		.Y(n_1170));

	NAND2X1 i_866(
		.A(acc[27]),
		.B(n_6195),
		.Y(n_1172));

	OAI21XL i_863(
		.A0(n_452),
		.A1(n_1172),
		.B0(n_863),
		.Y(n_1173));

	AOI31X1 i_864(
		.A0(n_6195),
		.A1(acc[29]),
		.A2(n_1031),
		.B0(n_1173),
		.Y(n_1174));

	OAI222XL i_862(
		.A0(n_548),
		.A1(n_1086),
		.B0(n_1152),
		.B1(n_4506),
		.C0(n_542),
		.C1(n_6306),
		.Y(n_1176));

	AOI222X1 i_859(
		.A0(ar1[14]),
		.A1(n_1026),
		.B0(acc[14]),
		.B1(n_4513),
		.C0(ar0[14]),
		.C1(n_1023),
		.Y(n_1179));

	AOI222XL i_857(
		.A0(p_data_out[14]),
		.A1(n_1035),
		.B0(port_data_out[14]),
		.B1(n_1015),
		.C0(mdr[14]),
		.C1(dmov_inc),
		.Y(n_1181));

	OAI222XL i_851(
		.A0(n_545),
		.A1(n_1086),
		.B0(n_452),
		.B1(n_1152),
		.C0(n_539),
		.C1(n_6306),
		.Y(n_1187));

	NAND4BXL i_854(
		.AN(n_1187),
		.B(n_851),
		.C(n_850),
		.D(n_852),
		.Y(n_1188));

	AOI222X1 i_848(
		.A0(ar1[15]),
		.A1(n_7152),
		.B0(acc[15]),
		.B1(n_4513),
		.C0(ar0[15]),
		.C1(n_7155),
		.Y(n_1190));

	AOI222X1 i_846(
		.A0(p_data_out[15]),
		.A1(n_7161),
		.B0(port_data_out[15]),
		.B1(n_7164),
		.C0(n_7112),
		.C1(mdr[15]),
		.Y(n_1192));

	MXI2X1 i_29(
		.S0(ir[7]),
		.B(ar[7]),
		.A(dp),
		.Y(n_1194));

	MXI2X1 i_578618(
		.S0(ir[7]),
		.B(ar[6]),
		.A(ir[6]),
		.Y(n_1195));

	MXI2X1 i_588619(
		.S0(ir[7]),
		.B(ar[5]),
		.A(ir[5]),
		.Y(n_1196));

	MXI2X1 i_24(
		.S0(ir[7]),
		.B(ar[4]),
		.A(ir[4]),
		.Y(n_1197));

	MXI2X1 i_608621(
		.S0(ir[7]),
		.B(ar_36576),
		.A(n_4524),
		.Y(n_1198));

	MXI2X1 i_18(
		.S0(ir[7]),
		.B(ar_26577),
		.A(n_4523),
		.Y(n_1199));

	MXI2X1 i_638624(
		.S0(ir[7]),
		.B(ar_06579),
		.A(n_4521),
		.Y(n_1200));

	MXI2X1 i_628623(
		.S0(ir[7]),
		.B(ar_16578),
		.A(n_4522),
		.Y(n_1201));

	NAND4X1 i_35(
		.A(n_1199),
		.B(dmov_inc),
		.C(n_1201),
		.D(n_1200),
		.Y(n_1204));

	NOR2BX1 i_59(
		.AN(n_1198),
		.B(n_1204),
		.Y(n_1205));

	NOR2BX1 i_17(
		.AN(n_1205),
		.B(n_1197),
		.Y(n_1206));

	NOR2BX1 i_54(
		.AN(n_1206),
		.B(n_1196),
		.Y(n_1207));

	NOR2BX1 i_67(
		.AN(n_1207),
		.B(n_1195),
		.Y(n_1208));

	NAND2X1 i_55(
		.A(dmov_inc),
		.B(n_1200),
		.Y(n_1209));

	NAND3X1 i_68(
		.A(dmov_inc),
		.B(n_1200),
		.C(n_1201),
		.Y(n_1210));

	NOR2X1 i_56(
		.A(sel_op_b[2]),
		.B(sel_op_b[0]),
		.Y(n_1211));

	NOR3BX1 i_2(
		.AN(sel_op_b[2]),
		.B(sel_op_b[0]),
		.C(sel_op_b[1]),
		.Y(n_1213));

	NOR2BX1 i_841(
		.AN(sel_op_b[0]),
		.B(sel_op_b[1]),
		.Y(n_1214));

	NOR2BX1 i_12(
		.AN(n_1214),
		.B(sel_op_b[2]),
		.Y(n_1215));

	AOI22X1 i_840(
		.A0(mdr[14]),
		.A1(n_7003),
		.B0(mdr[15]),
		.B1(n_1211),
		.Y(n_1216));

	NAND2X1 i_5(
		.A(ir[11]),
		.B(n_1211),
		.Y(n_1217));

	NAND3X1 i_28(
		.A(ir[11]),
		.B(n_1211),
		.C(port_addrs_in[2]),
		.Y(n_1218));

	AOI22X1 i_839(
		.A0(mdr[13]),
		.A1(n_7003),
		.B0(n_4496),
		.B1(n_4511),
		.Y(n_1219));

	NOR3X1 i_3(
		.A(sel_op_b[2]),
		.B(sel_op_b[0]),
		.C(ir[11]),
		.Y(n_1220));

	NAND2BX1 i_15(
		.AN(port_addrs_in[2]),
		.B(mdr[15]),
		.Y(n_1221));

	OAI21XL i_52(
		.A0(n_1217),
		.A1(n_1221),
		.B0(n_807),
		.Y(n_1222));

	AOI21X1 i_838(
		.A0(p[29]),
		.A1(n_7236),
		.B0(n_1222),
		.Y(n_1223));

	AOI21X1 i_835(
		.A0(p[28]),
		.A1(n_7236),
		.B0(n_1222),
		.Y(n_1226));

	AOI22X1 i_834(
		.A0(mdr[15]),
		.A1(n_7170),
		.B0(mdr[14]),
		.B1(n_7158),
		.Y(n_1227));

	AOI22X1 i_833(
		.A0(mdr[12]),
		.A1(n_4508),
		.B0(mdr[13]),
		.B1(n_7056),
		.Y(n_1228));

	AOI22X1 i_832(
		.A0(mdr[11]),
		.A1(n_7003),
		.B0(n_446),
		.B1(n_4511),
		.Y(n_1229));

	AOI21X1 i_831(
		.A0(p[27]),
		.A1(n_7236),
		.B0(n_1222),
		.Y(n_1230));

	AOI22X1 i_830(
		.A0(mdr[14]),
		.A1(n_7170),
		.B0(mdr[13]),
		.B1(n_7158),
		.Y(n_1231));

	AOI22X1 i_829(
		.A0(mdr[11]),
		.A1(n_4508),
		.B0(mdr[12]),
		.B1(n_7056),
		.Y(n_1232));

	AOI22X1 i_828(
		.A0(mdr[10]),
		.A1(n_7003),
		.B0(n_445),
		.B1(n_4511),
		.Y(n_1233));

	AOI21X1 i_827(
		.A0(p[26]),
		.A1(n_7236),
		.B0(n_1222),
		.Y(n_1234));

	AOI22X1 i_826(
		.A0(mdr[13]),
		.A1(n_7170),
		.B0(mdr[12]),
		.B1(n_7158),
		.Y(n_1235));

	AOI22X1 i_825(
		.A0(mdr[10]),
		.A1(n_4508),
		.B0(mdr[11]),
		.B1(n_7056),
		.Y(n_1236));

	NOR2X1 i_25(
		.A(port_addrs_in[2]),
		.B(n_1217),
		.Y(n_1237));

	AOI222X1 i_824(
		.A0(n_7001),
		.A1(n_4496),
		.B0(n_444),
		.B1(n_4511),
		.C0(mdr[9]),
		.C1(n_7003),
		.Y(n_1239));

	AOI22X1 i_821(
		.A0(mdr[12]),
		.A1(n_7170),
		.B0(mdr[11]),
		.B1(n_7158),
		.Y(n_1241));

	OAI22X1 i_818(
		.A0(n_447),
		.A1(n_4509),
		.B0(n_443),
		.B1(n_1218),
		.Y(n_1243));

	AOI21X1 i_819(
		.A0(mdr[8]),
		.A1(n_7003),
		.B0(n_1243),
		.Y(n_1244));

	AOI22X1 i_816(
		.A0(mdr[11]),
		.A1(n_7170),
		.B0(mdr[10]),
		.B1(n_7158),
		.Y(n_1246));

	AOI22X1 i_815(
		.A0(mdr[8]),
		.A1(n_4508),
		.B0(mdr[9]),
		.B1(n_7056),
		.Y(n_1247));

	AOI222X1 i_814(
		.A0(n_446),
		.A1(n_7001),
		.B0(n_442),
		.B1(n_4511),
		.C0(mdr[7]),
		.C1(n_7003),
		.Y(n_1249));

	AOI22X1 i_811(
		.A0(mdr[10]),
		.A1(n_7170),
		.B0(mdr[9]),
		.B1(n_7158),
		.Y(n_1251));

	AOI22X1 i_810(
		.A0(mdr[7]),
		.A1(n_4508),
		.B0(mdr[8]),
		.B1(n_7056),
		.Y(n_1252));

	AOI222X1 i_809(
		.A0(n_445),
		.A1(n_7001),
		.B0(n_441),
		.B1(n_4511),
		.C0(mdr[6]),
		.C1(n_7003),
		.Y(n_1254));

	AOI22X1 i_806(
		.A0(mdr[9]),
		.A1(n_7170),
		.B0(mdr[8]),
		.B1(n_7158),
		.Y(n_1256));

	AOI22X1 i_805(
		.A0(mdr[6]),
		.A1(n_4508),
		.B0(mdr[7]),
		.B1(n_7056),
		.Y(n_1257));

	NAND2X1 i_26(
		.A(port_addrs_in[2]),
		.B(n_1220),
		.Y(n_1258));

	AOI222X1 i_804(
		.A0(n_4496),
		.A1(n_4507),
		.B0(n_440),
		.B1(n_4511),
		.C0(n_444),
		.C1(n_7001),
		.Y(n_1260));

	AOI22X1 i_801(
		.A0(p[21]),
		.A1(n_7236),
		.B0(mdr[5]),
		.B1(n_7003),
		.Y(n_1261));

	AOI22X1 i_800(
		.A0(mdr[8]),
		.A1(n_7170),
		.B0(mdr[7]),
		.B1(n_7158),
		.Y(n_1263));

	AOI22X1 i_799(
		.A0(mdr[5]),
		.A1(n_4508),
		.B0(mdr[6]),
		.B1(n_7056),
		.Y(n_1264));

	OAI222XL i_798(
		.A0(n_447),
		.A1(n_1258),
		.B0(n_1218),
		.B1(n_4498),
		.C0(n_443),
		.C1(n_4509),
		.Y(n_1266));

	AOI22X1 i_795(
		.A0(p[20]),
		.A1(n_7236),
		.B0(mdr[4]),
		.B1(n_7003),
		.Y(n_1267));

	AOI22X1 i_794(
		.A0(mdr[7]),
		.A1(n_7170),
		.B0(mdr[6]),
		.B1(n_7158),
		.Y(n_1269));

	AOI22X1 i_793(
		.A0(mdr[4]),
		.A1(n_4508),
		.B0(mdr[5]),
		.B1(n_7056),
		.Y(n_1270));

	AOI211X1 i_792(
		.A0(n_442),
		.A1(n_7001),
		.B0(n_758),
		.C0(n_757),
		.Y(n_1272));

	AOI22X1 i_789(
		.A0(p[19]),
		.A1(n_7236),
		.B0(mdr[3]),
		.B1(n_7003),
		.Y(n_1273));

	AOI22X1 i_788(
		.A0(mdr[6]),
		.A1(n_7170),
		.B0(mdr[5]),
		.B1(n_7158),
		.Y(n_1275));

	AOI22X1 i_787(
		.A0(mdr[3]),
		.A1(n_4508),
		.B0(mdr[4]),
		.B1(n_7056),
		.Y(n_1276));

	AOI222X1 i_786(
		.A0(n_445),
		.A1(n_4507),
		.B0(n_437),
		.B1(n_4511),
		.C0(n_441),
		.C1(n_7001),
		.Y(n_1278));

	AOI22X1 i_783(
		.A0(p[18]),
		.A1(n_1213),
		.B0(mdr[2]),
		.B1(n_7003),
		.Y(n_1279));

	AOI22X1 i_782(
		.A0(mdr[5]),
		.A1(n_7170),
		.B0(mdr[4]),
		.B1(n_7158),
		.Y(n_1281));

	AOI22X1 i_781(
		.A0(mdr[2]),
		.A1(n_4508),
		.B0(mdr[3]),
		.B1(n_7056),
		.Y(n_1282));

	NAND2BX1 i_27(
		.AN(port_addrs_in[2]),
		.B(n_1220),
		.Y(n_1283));

	OAI222XL i_780(
		.A0(n_1283),
		.A1(n_449),
		.B0(n_4499),
		.B1(n_1218),
		.C0(n_1258),
		.C1(n_4497),
		.Y(n_1285));

	AOI222X1 i_778(
		.A0(mdr[1]),
		.A1(n_7003),
		.B0(n_440),
		.B1(n_7001),
		.C0(p[17]),
		.C1(n_7236),
		.Y(n_1287));

	AOI22X1 i_776(
		.A0(mdr[4]),
		.A1(n_7170),
		.B0(mdr[3]),
		.B1(n_7158),
		.Y(n_1288));

	AOI22X1 i_775(
		.A0(mdr[1]),
		.A1(n_4508),
		.B0(mdr[2]),
		.B1(n_7056),
		.Y(n_1289));

	OAI222XL i_774(
		.A0(n_447),
		.A1(n_1283),
		.B0(n_1218),
		.B1(n_4500),
		.C0(n_1258),
		.C1(n_443),
		.Y(n_1291));

	AOI222X1 i_772(
		.A0(mdr[0]),
		.A1(n_7003),
		.B0(n_7001),
		.B1(n_439),
		.C0(p[16]),
		.C1(n_7236),
		.Y(n_1293));

	AOI22X1 i_770(
		.A0(mdr[3]),
		.A1(n_7170),
		.B0(mdr[2]),
		.B1(n_7158),
		.Y(n_1294));

	AOI22X1 i_767(
		.A0(n_446),
		.A1(n_4505),
		.B0(n_4511),
		.B1(n_430),
		.Y(n_1295));

	AOI22X1 i_766(
		.A0(n_438),
		.A1(n_7001),
		.B0(n_442),
		.B1(n_4507),
		.Y(n_1296));

	NAND2X1 i_11(
		.A(sel_op_b[2]),
		.B(n_1214),
		.Y(n_1298));

	NOR2BX1 i_10(
		.AN(sel_op_b[1]),
		.B(n_1211),
		.Y(n_1299));

	AOI22X1 i_764(
		.A0(p[15]),
		.A1(n_7006),
		.B0(mdr[15]),
		.B1(n_7247),
		.Y(n_1300));

	AOI22X1 i_761(
		.A0(n_445),
		.A1(n_4505),
		.B0(n_4511),
		.B1(n_4502),
		.Y(n_1303));

	AOI22X1 i_760(
		.A0(n_437),
		.A1(n_7001),
		.B0(n_441),
		.B1(n_4507),
		.Y(n_1304));

	AOI22X1 i_758(
		.A0(p[14]),
		.A1(n_1213),
		.B0(mdr[14]),
		.B1(n_7247),
		.Y(n_1306));

	NOR2X1 i_64(
		.A(n_432),
		.B(port_addrs_in[1]),
		.Y(n_1308));

	AOI22X1 i_756(
		.A0(n_444),
		.A1(n_4505),
		.B0(n_1308),
		.B1(n_4511),
		.Y(n_1309));

	AOI22X1 i_755(
		.A0(n_7001),
		.A1(n_436),
		.B0(n_440),
		.B1(n_4507),
		.Y(n_1310));

	AOI22X1 i_753(
		.A0(p[13]),
		.A1(n_7006),
		.B0(mdr[13]),
		.B1(n_7247),
		.Y(n_1312));

	NAND2X1 i_34(
		.A(mdr[0]),
		.B(n_7170),
		.Y(n_1314));

	AOI2BB1X1 i_751(
		.A0N(n_443),
		.A1N(n_1283),
		.B0(n_701),
		.Y(n_1315));

	AOI22X1 i_750(
		.A0(n_435),
		.A1(n_7001),
		.B0(n_439),
		.B1(n_4507),
		.Y(n_1316));

	AOI22X1 i_748(
		.A0(p[12]),
		.A1(n_7006),
		.B0(mdr[12]),
		.B1(n_7247),
		.Y(n_1318));

	AOI22X1 i_746(
		.A0(n_438),
		.A1(n_4507),
		.B0(n_442),
		.B1(n_4505),
		.Y(n_1320));

	AOI222X1 i_745(
		.A0(mdr[11]),
		.A1(n_7247),
		.B0(ir[11]),
		.B1(n_4504),
		.C0(p[11]),
		.C1(n_7006),
		.Y(n_1323));

	AOI22X1 i_742(
		.A0(n_437),
		.A1(n_4507),
		.B0(n_441),
		.B1(n_4505),
		.Y(n_1324));

	AOI222X1 i_741(
		.A0(mdr[10]),
		.A1(n_7247),
		.B0(port_addrs_in[2]),
		.B1(n_4504),
		.C0(p[10]),
		.C1(n_7006),
		.Y(n_1327));

	AOI22X1 i_738(
		.A0(n_440),
		.A1(n_4505),
		.B0(n_1308),
		.B1(n_7001),
		.Y(n_1328));

	AOI222X1 i_737(
		.A0(mdr[9]),
		.A1(n_7247),
		.B0(port_addrs_in[1]),
		.B1(n_4504),
		.C0(p[9]),
		.C1(n_7006),
		.Y(n_1331));

	AOI22X1 i_734(
		.A0(n_4507),
		.A1(n_435),
		.B0(n_439),
		.B1(n_4505),
		.Y(n_1332));

	AOI222X1 i_733(
		.A0(mdr[8]),
		.A1(n_7247),
		.B0(port_addrs_in[0]),
		.B1(n_4504),
		.C0(p[8]),
		.C1(n_7006),
		.Y(n_1335));

	AOI22X1 i_730(
		.A0(n_430),
		.A1(n_4507),
		.B0(n_438),
		.B1(n_4505),
		.Y(n_1336));

	AOI22X1 i_729(
		.A0(p[7]),
		.A1(n_7006),
		.B0(mdr[7]),
		.B1(n_7247),
		.Y(n_1338));

	AOI22X1 i_727(
		.A0(n_4502),
		.A1(n_4507),
		.B0(n_437),
		.B1(n_4505),
		.Y(n_1339));

	AOI22X1 i_726(
		.A0(p[6]),
		.A1(n_7006),
		.B0(mdr[6]),
		.B1(n_1299),
		.Y(n_1341));

	OAI21XL i_724(
		.A0(n_4499),
		.A1(n_1283),
		.B0(n_660),
		.Y(n_1342));

	AOI31X1 i_725(
		.A0(sel_op_b[2]),
		.A1(ir[5]),
		.A2(n_1214),
		.B0(n_1342),
		.Y(n_1343));

	AOI22X1 i_723(
		.A0(p[5]),
		.A1(n_7006),
		.B0(mdr[5]),
		.B1(n_7247),
		.Y(n_1344));

	AOI32X1 i_721(
		.A0(mdr[0]),
		.A1(n_7170),
		.A2(n_4507),
		.B0(n_435),
		.B1(n_4505),
		.Y(n_1345));

	AOI22X1 i_720(
		.A0(p[4]),
		.A1(n_7006),
		.B0(mdr[4]),
		.B1(n_7247),
		.Y(n_1347));

	AOI22X1 i_718(
		.A0(p[3]),
		.A1(n_7006),
		.B0(mdr[3]),
		.B1(n_7247),
		.Y(n_1349));

	AOI22X1 i_716(
		.A0(p[2]),
		.A1(n_7006),
		.B0(mdr[2]),
		.B1(n_1299),
		.Y(n_1351));

	AOI32X1 i_715(
		.A0(sel_op_b[2]),
		.A1(n_1214),
		.A2(ir[1]),
		.B0(n_1308),
		.B1(n_4505),
		.Y(n_1352));

	AOI22X1 i_714(
		.A0(p[1]),
		.A1(n_7006),
		.B0(mdr[1]),
		.B1(n_1299),
		.Y(n_1353));

	AOI22X1 i_712(
		.A0(p[0]),
		.A1(n_7006),
		.B0(mdr[0]),
		.B1(n_1299),
		.Y(n_1355));

	NOR3BX1 i_1(
		.AN(sel_op_a[0]),
		.B(sel_op_a[1]),
		.C(sel_op_a[2]),
		.Y(n_1357));

	NAND2X1 i_710(
		.A(sel_op_a[1]),
		.B(sel_op_a[0]),
		.Y(n_1358));

	NOR2X1 i_8(
		.A(n_1358),
		.B(sel_op_a[2]),
		.Y(n_1359));

	AOI22X1 i_709(
		.A0(acc[15]),
		.A1(n_7015),
		.B0(top[15]),
		.B1(n_7239),
		.Y(n_1360));

	AOI22X1 i_708(
		.A0(acc[14]),
		.A1(n_1357),
		.B0(top[14]),
		.B1(n_7239),
		.Y(n_1361));

	AOI22X1 i_707(
		.A0(acc[13]),
		.A1(n_7015),
		.B0(top[13]),
		.B1(n_7239),
		.Y(n_1362));

	AOI22X1 i_706(
		.A0(acc[12]),
		.A1(n_7015),
		.B0(top[12]),
		.B1(n_7239),
		.Y(n_1363));

	AOI22X1 i_705(
		.A0(acc[11]),
		.A1(n_7015),
		.B0(top[11]),
		.B1(n_7239),
		.Y(n_1364));

	AOI22X1 i_704(
		.A0(acc[10]),
		.A1(n_7015),
		.B0(top[10]),
		.B1(n_7239),
		.Y(n_1365));

	AOI22X1 i_703(
		.A0(acc[9]),
		.A1(n_7015),
		.B0(top[9]),
		.B1(n_7239),
		.Y(n_1366));

	AOI22X1 i_702(
		.A0(acc[8]),
		.A1(n_7015),
		.B0(top[8]),
		.B1(n_7239),
		.Y(n_1367));

	NOR2X1 i_14(
		.A(n_1358),
		.B(n_4520),
		.Y(n_1368));

	AOI22X1 i_700(
		.A0(top[7]),
		.A1(n_7239),
		.B0(ir[7]),
		.B1(n_1368),
		.Y(n_1369));

	AOI22X1 i_699(
		.A0(mdr[7]),
		.A1(n_7227),
		.B0(acc[7]),
		.B1(n_7015),
		.Y(n_1370));

	AOI22X1 i_698(
		.A0(top[6]),
		.A1(n_1359),
		.B0(ir[6]),
		.B1(n_1368),
		.Y(n_1371));

	AOI22X1 i_697(
		.A0(mdr[6]),
		.A1(n_410),
		.B0(acc[6]),
		.B1(n_7015),
		.Y(n_1372));

	AOI22X1 i_696(
		.A0(top[5]),
		.A1(n_7239),
		.B0(ir[5]),
		.B1(n_1368),
		.Y(n_1373));

	AOI22X1 i_695(
		.A0(mdr[5]),
		.A1(n_7227),
		.B0(acc[5]),
		.B1(n_7015),
		.Y(n_1374));

	AOI22X1 i_694(
		.A0(top[4]),
		.A1(n_1359),
		.B0(ir[4]),
		.B1(n_1368),
		.Y(n_1375));

	AOI22X1 i_693(
		.A0(mdr[4]),
		.A1(n_7227),
		.B0(acc[4]),
		.B1(n_7015),
		.Y(n_1376));

	AOI22X1 i_691(
		.A0(mdr[3]),
		.A1(n_7227),
		.B0(acc[3]),
		.B1(n_7015),
		.Y(n_1378));

	AOI22X1 i_689(
		.A0(mdr[2]),
		.A1(n_7227),
		.B0(acc[2]),
		.B1(n_7015),
		.Y(n_1380));

	AOI22X1 i_688(
		.A0(top[1]),
		.A1(n_1359),
		.B0(ir[1]),
		.B1(n_1368),
		.Y(n_1381));

	AOI22X1 i_687(
		.A0(mdr[1]),
		.A1(n_410),
		.B0(n_7015),
		.B1(acc[1]),
		.Y(n_1382));

	AOI22X1 i_685(
		.A0(mdr[0]),
		.A1(n_7227),
		.B0(n_7015),
		.B1(acc[0]),
		.Y(n_1384));

	OR2X1 i_5354(
		.A(enc_go_prog),
		.B(dec_go_prog),
		.Y(go_prog));

	OR2X1 i_5356(
		.A(enc_go_port),
		.B(dec_go_port),
		.Y(go_port));

	OR2X1 i_5357(
		.A(enc_go_data),
		.B(dec_go_data),
		.Y(go_data));

	OR2X1 i_5358(
		.A(enc_read_data),
		.B(dec_read_data),
		.Y(read_data));

	OR2X1 i_5366(
		.A(enc_read_prog),
		.B(dec_read_prog),
		.Y(read_prog));

	OR2X1 i_5369(
		.A(enc_read_port),
		.B(dec_read_port),
		.Y(read_port));

	NAND4BXL i_5427(
		.AN(n_1052),
		.B(n_1056),
		.C(n_1055),
		.D(n_1044),
		.Y(data_in[0]));

	NAND4BXL i_5434(
		.AN(n_1061),
		.B(n_1065),
		.C(n_1064),
		.D(n_1059),
		.Y(data_in[1]));

	NAND4BXL i_5441(
		.AN(n_1068),
		.B(n_1075),
		.C(n_1074),
		.D(n_1071),
		.Y(data_in[2]));

	NAND4BXL i_5448(
		.AN(n_1078),
		.B(n_1084),
		.C(n_1083),
		.D(n_1080),
		.Y(data_in[3]));

	NAND4BXL i_5455(
		.AN(n_1088),
		.B(n_1093),
		.C(n_1092),
		.D(n_1089),
		.Y(data_in[4]));

	NAND4BXL i_5462(
		.AN(n_1096),
		.B(n_1101),
		.C(n_1100),
		.D(n_1097),
		.Y(data_in[5]));

	NAND4BXL i_5469(
		.AN(n_1104),
		.B(n_1109),
		.C(n_1108),
		.D(n_1105),
		.Y(data_in[6]));

	NAND4BXL i_5476(
		.AN(n_1112),
		.B(n_1117),
		.C(n_1116),
		.D(n_1113),
		.Y(data_in[7]));

	NAND4BXL i_5483(
		.AN(n_1120),
		.B(n_1125),
		.C(n_1124),
		.D(n_1121),
		.Y(data_in[8]));

	NAND4BXL i_5490(
		.AN(n_1128),
		.B(n_1133),
		.C(n_1132),
		.D(n_1129),
		.Y(data_in[9]));

	NAND4BXL i_5497(
		.AN(n_1136),
		.B(n_1141),
		.C(n_1140),
		.D(n_1137),
		.Y(data_in[10]));

	NAND4BXL i_5504(
		.AN(n_1144),
		.B(n_1149),
		.C(n_1148),
		.D(n_1145),
		.Y(data_in[11]));

	NAND4BXL i_5511(
		.AN(n_1154),
		.B(n_1160),
		.C(n_1159),
		.D(n_1156),
		.Y(data_in[12]));

	NAND4BXL i_5518(
		.AN(n_1164),
		.B(n_1170),
		.C(n_1169),
		.D(n_1166),
		.Y(data_in[13]));

	NAND4BXL i_5525(
		.AN(n_1176),
		.B(n_1181),
		.C(n_1179),
		.D(n_1174),
		.Y(data_in[14]));

	NAND3BX1 i_5532(
		.AN(n_1188),
		.B(n_1192),
		.C(n_1190),
		.Y(data_in[15]));

	MX2X1 i_248287(
		.S0(n_6255),
		.B(ar1[15]),
		.A(ar0[15]),
		.Y(ar[15]));

	MX2X1 i_258288(
		.S0(n_6255),
		.B(ar1[14]),
		.A(ar0[14]),
		.Y(ar[14]));

	MX2X1 i_268289(
		.S0(n_6255),
		.B(ar1[13]),
		.A(ar0[13]),
		.Y(ar[13]));

	MX2X1 i_278290(
		.S0(n_6255),
		.B(ar1[12]),
		.A(ar0[12]),
		.Y(ar[12]));

	MX2X1 i_288291(
		.S0(n_6255),
		.B(ar1[11]),
		.A(ar0[11]),
		.Y(ar[11]));

	MX2X1 i_298292(
		.S0(n_6255),
		.B(ar1[10]),
		.A(ar0[10]),
		.Y(ar[10]));

	MX2X1 i_308293(
		.S0(n_6255),
		.B(ar1[9]),
		.A(ar0[9]),
		.Y(ar[9]));

	MX2X1 i_318294(
		.S0(n_6255),
		.B(ar1[8]),
		.A(ar0[8]),
		.Y(ar[8]));

	MX2X1 i_328295(
		.S0(n_6255),
		.B(ar1[7]),
		.A(ar0[7]),
		.Y(ar[7]));

	MX2X1 i_338296(
		.S0(n_6255),
		.B(ar1[6]),
		.A(ar0[6]),
		.Y(ar[6]));

	MX2X1 i_348297(
		.S0(n_6255),
		.B(ar1[5]),
		.A(ar0[5]),
		.Y(ar[5]));

	MX2X1 i_358298(
		.S0(n_7084),
		.B(ar1[4]),
		.A(ar0[4]),
		.Y(ar[4]));

	MXI2X1 i_368299(
		.S0(n_7084),
		.B(ar1[3]),
		.A(ar0[3]),
		.Y(ar_36576));

	MXI2X1 i_378300(
		.S0(n_7084),
		.B(ar1[2]),
		.A(ar0[2]),
		.Y(ar_26577));

	MXI2X1 i_388301(
		.S0(n_7084),
		.B(ar1[1]),
		.A(ar0[1]),
		.Y(ar_16578));

	MXI2X1 i_398302(
		.S0(n_7084),
		.B(ar1[0]),
		.A(ar0[0]),
		.Y(ar_06579));

	OAI21XL i_568625(
		.A0(n_1208),
		.A1(n_1194),
		.B0(n_489),
		.Y(addrs_in[7]));

	OAI21XL i_578626(
		.A0(n_1207),
		.A1(n_1195),
		.B0(n_487),
		.Y(addrs_in[6]));

	OAI21XL i_588627(
		.A0(n_1206),
		.A1(n_1196),
		.B0(n_485),
		.Y(addrs_in[5]));

	OAI21XL i_598628(
		.A0(n_1205),
		.A1(n_1197),
		.B0(n_483),
		.Y(addrs_in[4]));

	OAI21XL i_608629(
		.A0(n_1204),
		.A1(n_1198),
		.B0(n_482),
		.Y(addrs_in[3]));

	OAI21XL i_618630(
		.A0(n_1210),
		.A1(n_1199),
		.B0(n_480),
		.Y(addrs_in[2]));

	OAI21XL i_628631(
		.A0(n_1209),
		.A1(n_1201),
		.B0(n_478),
		.Y(addrs_in[1]));

	XOR2X1 i_638632(
		.A(n_1200),
		.B(dmov_inc),
		.Y(addrs_in[0]));

	MX2X1 i_582(
		.S0(pc_acc),
		.B(acc[7]),
		.A(pc[7]),
		.Y(p_addrs_in[7]));

	MX2X1 i_583(
		.S0(pc_acc),
		.B(acc[6]),
		.A(pc[6]),
		.Y(p_addrs_in[6]));

	MX2X1 i_584(
		.S0(pc_acc),
		.B(acc[5]),
		.A(pc[5]),
		.Y(p_addrs_in[5]));

	MX2X1 i_585(
		.S0(pc_acc),
		.B(acc[4]),
		.A(pc[4]),
		.Y(p_addrs_in[4]));

	MX2X1 i_586(
		.S0(pc_acc),
		.B(acc[3]),
		.A(pc[3]),
		.Y(p_addrs_in[3]));

	MX2X1 i_587(
		.S0(pc_acc),
		.B(acc[2]),
		.A(pc[2]),
		.Y(p_addrs_in[2]));

	MX2X1 i_588(
		.S0(pc_acc),
		.B(acc[1]),
		.A(pc[1]),
		.Y(p_addrs_in[1]));

	MX2X1 i_589(
		.S0(pc_acc),
		.B(acc[0]),
		.A(pc[0]),
		.Y(p_addrs_in[0]));

	AOI22X1 i_517(
		.A0(p[31]),
		.A1(n_7236),
		.B0(mdr[15]),
		.B1(n_456),
		.Y(opb_316580));

	OAI2BB1X1 i_518(
		.A0N(p[30]),
		.A1N(n_7236),
		.B0(n_1216),
		.Y(opb[30]));

	NAND2X1 i_519(
		.A(n_1223),
		.B(n_1219),
		.Y(opb[29]));

	OAI211X1 i_520(
		.A0(n_447),
		.A1(n_1218),
		.B0(n_832),
		.C0(n_1226),
		.Y(opb[28]));

	NAND2X1 i_521(
		.A(n_1230),
		.B(n_1229),
		.Y(opb[27]));

	NAND2X1 i_522(
		.A(n_1234),
		.B(n_1233),
		.Y(opb[26]));

	NAND3X1 i_523(
		.A(n_808),
		.B(n_807),
		.C(n_1239),
		.Y(opb[25]));

	NAND3X1 i_524(
		.A(n_807),
		.B(n_799),
		.C(n_1244),
		.Y(opb[24]));

	NAND3X1 i_525(
		.A(n_807),
		.B(n_791),
		.C(n_1249),
		.Y(opb[23]));

	NAND3X1 i_526(
		.A(n_807),
		.B(n_783),
		.C(n_1254),
		.Y(opb[22]));

	NAND3X1 i_527(
		.A(n_775),
		.B(n_1261),
		.C(n_1260),
		.Y(opb[21]));

	NAND3X1 i_528(
		.A(n_775),
		.B(n_1267),
		.C(n_4512),
		.Y(opb[20]));

	NAND3X1 i_529(
		.A(n_775),
		.B(n_1273),
		.C(n_1272),
		.Y(opb[19]));

	NAND3X1 i_530(
		.A(n_775),
		.B(n_1279),
		.C(n_1278),
		.Y(opb[18]));

	NAND2BX1 i_531(
		.AN(n_1285),
		.B(n_1287),
		.Y(opb[17]));

	NAND2BX1 i_532(
		.AN(n_1291),
		.B(n_1293),
		.Y(opb[16]));

	NAND4X1 i_533(
		.A(n_719),
		.B(n_1300),
		.C(n_1296),
		.D(n_1295),
		.Y(opb[15]));

	NAND4X1 i_534(
		.A(n_719),
		.B(n_1306),
		.C(n_1304),
		.D(n_1303),
		.Y(opb[14]));

	NAND4X1 i_535(
		.A(n_719),
		.B(n_1312),
		.C(n_1310),
		.D(n_1309),
		.Y(opb[13]));

	NAND4X1 i_536(
		.A(n_719),
		.B(n_1318),
		.C(n_1316),
		.D(n_1315),
		.Y(opb[12]));

	OAI211X1 i_537(
		.A0(n_4501),
		.A1(n_4509),
		.B0(n_1320),
		.C0(n_1323),
		.Y(opb[11]));

	OAI211X1 i_538(
		.A0(n_428),
		.A1(n_4509),
		.B0(n_1324),
		.C0(n_1327),
		.Y(opb[10]));

	OAI211X1 i_539(
		.A0(n_1258),
		.A1(n_4499),
		.B0(n_1328),
		.C0(n_1331),
		.Y(opb[9]));

	OAI211X1 i_540(
		.A0(n_1314),
		.A1(n_4509),
		.B0(n_1332),
		.C0(n_1335),
		.Y(opb[8]));

	NAND3X1 i_541(
		.A(n_672),
		.B(n_1338),
		.C(n_1336),
		.Y(opb[7]));

	NAND3X1 i_542(
		.A(n_667),
		.B(n_1341),
		.C(n_1339),
		.Y(opb[6]));

	NAND2X1 i_543(
		.A(n_1344),
		.B(n_1343),
		.Y(opb[5]));

	NAND3X1 i_544(
		.A(n_657),
		.B(n_1347),
		.C(n_1345),
		.Y(opb[4]));

	OAI221XL i_545(
		.A0(n_1298),
		.A1(n_4524),
		.B0(n_4501),
		.B1(n_1283),
		.C0(n_1349),
		.Y(\nbus_686[3] ));

	OAI221XL i_546(
		.A0(n_1298),
		.A1(n_4523),
		.B0(n_428),
		.B1(n_1283),
		.C0(n_1351),
		.Y(\nbus_684[2] ));

	NAND2X1 i_547(
		.A(n_1353),
		.B(n_1352),
		.Y(opb[1]));

	OAI221XL i_548(
		.A0(n_1298),
		.A1(n_4521),
		.B0(n_1314),
		.B1(n_1283),
		.C0(n_1355),
		.Y(\nbus_683[0] ));

	OAI2BB1X1 i_5178960(
		.A0N(acc[31]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[31]));

	OAI2BB1X1 i_5188961(
		.A0N(acc[30]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[30]));

	OAI2BB1X1 i_5198962(
		.A0N(acc[29]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[29]));

	OAI2BB1X1 i_5208963(
		.A0N(acc[28]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[28]));

	OAI2BB1X1 i_5218964(
		.A0N(acc[27]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[27]));

	OAI2BB1X1 i_5228965(
		.A0N(acc[26]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[26]));

	OAI2BB1X1 i_5238966(
		.A0N(acc[25]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[25]));

	OAI2BB1X1 i_5248967(
		.A0N(acc[24]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[24]));

	OAI2BB1X1 i_5258968(
		.A0N(acc[23]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[23]));

	OAI2BB1X1 i_5268969(
		.A0N(acc[22]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[22]));

	OAI2BB1X1 i_5278970(
		.A0N(acc[21]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[21]));

	OAI2BB1X1 i_5288971(
		.A0N(acc[20]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[20]));

	OAI2BB1X1 i_5298972(
		.A0N(acc[19]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[19]));

	OAI2BB1X1 i_5308973(
		.A0N(acc[18]),
		.A1N(n_1357),
		.B0(n_402),
		.Y(opa[18]));

	OAI2BB1X1 i_5318974(
		.A0N(acc[17]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[17]));

	OAI2BB1X1 i_5328975(
		.A0N(acc[16]),
		.A1N(n_7224),
		.B0(n_7230),
		.Y(opa[16]));

	NAND2X1 i_5338976(
		.A(n_402),
		.B(n_1360),
		.Y(opa[15]));

	OAI2BB1X1 i_5348977(
		.A0N(mdr[14]),
		.A1N(n_7227),
		.B0(n_1361),
		.Y(opa[14]));

	OAI2BB1X1 i_5358978(
		.A0N(mdr[13]),
		.A1N(n_7227),
		.B0(n_1362),
		.Y(opa[13]));

	OAI2BB1X1 i_5368979(
		.A0N(mdr[12]),
		.A1N(n_7227),
		.B0(n_1363),
		.Y(opa[12]));

	OAI2BB1X1 i_5378980(
		.A0N(mdr[11]),
		.A1N(n_7227),
		.B0(n_1364),
		.Y(opa[11]));

	OAI2BB1X1 i_5388981(
		.A0N(mdr[10]),
		.A1N(n_7227),
		.B0(n_1365),
		.Y(opa[10]));

	OAI2BB1X1 i_5398982(
		.A0N(mdr[9]),
		.A1N(n_7227),
		.B0(n_1366),
		.Y(opa[9]));

	OAI2BB1X1 i_5408983(
		.A0N(mdr[8]),
		.A1N(n_7227),
		.B0(n_1367),
		.Y(opa[8]));

	NAND2X1 i_5418984(
		.A(n_1370),
		.B(n_1369),
		.Y(opa[7]));

	NAND2X1 i_5428985(
		.A(n_1372),
		.B(n_1371),
		.Y(opa[6]));

	NAND2X1 i_5438986(
		.A(n_1374),
		.B(n_1373),
		.Y(opa[5]));

	NAND2X1 i_5448987(
		.A(n_1376),
		.B(n_1375),
		.Y(opa[4]));

	OAI211X1 i_5458988(
		.A0(n_4503),
		.A1(n_4524),
		.B0(n_604),
		.C0(n_1378),
		.Y(opa[3]));

	OAI211X1 i_5468989(
		.A0(n_4503),
		.A1(n_4523),
		.B0(n_600),
		.C0(n_1380),
		.Y(\nbus_685[2] ));

	NAND2X1 i_5478990(
		.A(n_1382),
		.B(n_1381),
		.Y(opa[1]));

	OAI211X1 i_5488991(
		.A0(n_4503),
		.A1(n_4521),
		.B0(n_592),
		.C0(n_1384),
		.Y(opa[0]));

	INVX1 i_6102(
		.A(n_449),
		.Y(n_4496));

	INVX1 i_6103(
		.A(n_444),
		.Y(n_4497));

	INVX1 i_6104(
		.A(n_439),
		.Y(n_4498));

	INVX1 i_6105(
		.A(n_436),
		.Y(n_4499));

	INVX1 i_6106(
		.A(n_435),
		.Y(n_4500));

	INVX1 i_6107(
		.A(n_430),
		.Y(n_4501));

	INVX1 i_6108(
		.A(n_428),
		.Y(n_4502));

	INVX1 i_6109(
		.A(n_1368),
		.Y(n_4503));

	INVX1 i_6110(
		.A(n_1298),
		.Y(n_4504));

	INVX1 i_6111(
		.A(n_1283),
		.Y(n_4505));

	INVX1 i_6112(
		.A(n_7056),
		.Y(n_4506));

	INVX1 i_6113(
		.A(n_1258),
		.Y(n_4507));

	INVX1 i_6114(
		.A(n_452),
		.Y(n_4508));

	INVX1 i_6115(
		.A(n_7001),
		.Y(n_4509));

	INVX1 i_6116(
		.A(n_1241),
		.Y(n_4510));

	INVX1 i_6117(
		.A(n_1218),
		.Y(n_4511));

	INVX1 i_6118(
		.A(n_1266),
		.Y(n_4512));

	INVX1 i_6119(
		.A(n_1046),
		.Y(n_4513));

	INVX1 i_6120(
		.A(n_1152),
		.Y(n_4514));

	INVX1 i_6121(
		.A(opb_316580),
		.Y(opb[31]));

	INVX1 i_6122(
		.A(ar_06579),
		.Y(ar[0]));

	INVX1 i_6123(
		.A(ar_16578),
		.Y(ar[1]));

	INVX1 i_6124(
		.A(ar_26577),
		.Y(ar[2]));

	INVX1 i_6125(
		.A(ar_36576),
		.Y(ar[3]));

	INVX1 i_6126(
		.A(sel_op_a[2]),
		.Y(n_4520));

	INVX1 i_6127(
		.A(ir[0]),
		.Y(n_4521));

	INVX1 i_6128(
		.A(ir[1]),
		.Y(n_4522));

	INVX1 i_6129(
		.A(ir[2]),
		.Y(n_4523));

	INVX1 i_6130(
		.A(ir[3]),
		.Y(n_4524));

	INVX1 i_6131(
		.A(port_addrs_in[1]),
		.Y(n_4525));

	INVX1 i_6132(
		.A(acc[0]),
		.Y(n_4526));

	INVX1 i_6133(
		.A(acc[1]),
		.Y(n_4527));

endmodule
module tdsp_core_mach(
		samp_bio,
		samp_int,
		phi_1,
		phi_2,
		phi_3,
		phi_4,
		phi_5,
		phi_6,
		reset,
		clk,
		bus_request,
		bus_grant,
		bio,
		int,
		scan_en,
		BG_scan_in,
		BG_scan_out,
	FE_PT1_,
	SPCASCAN_N31_tdsp_state_2_,
	SPCASCAN_N32_two_cycle,
	FE_PT2_,
	SPCASCAN_N33_samp_int,
	SPCASCAN_N34_two_cycle,
	SPCASCAN_N35_three_cycle,
	FE_PT3_,
	SPCASCAN_N36_tdsp_state_1_,
	FE_PT4_);
   input FE_PT1_;
   output SPCASCAN_N31_tdsp_state_2_;
   input SPCASCAN_N32_two_cycle;
   input FE_PT2_;
   output SPCASCAN_N33_samp_int;
   input SPCASCAN_N34_two_cycle;
   input SPCASCAN_N35_three_cycle;
   input FE_PT3_;
   output SPCASCAN_N36_tdsp_state_1_;
   input FE_PT4_;

	output samp_bio;
	output samp_int;
	output phi_1;
	output phi_2;
	output phi_3;
	output phi_4;
	output phi_5;
	output phi_6;
	input reset;
	input clk;
	input bus_request;
	input bus_grant;
	input bio;
	input int;
	input scan_en;
	input BG_scan_in;
	output BG_scan_out;

	wire [2:0] tdsp_state;



	CLKBUFXL i_10014(
		.A(BG_scan_out),
		.Y(phi_6));

	NAND2X1 i_12(
		.A(n_102),
		.B(n_47),
		.Y(n_27));

	NAND4BXL i_122(
		.AN(n_45),
		.B(n_72),
		.C(n_22),
		.D(n_23),
		.Y(n_24));

	NAND2X1 i_14(
		.A(n_35),
		.B(n_2818),
		.Y(n_23));

	AOI32X1 i_228675(
		.A0(SPCASCAN_N31_tdsp_state_2_),
		.A1(SPCASCAN_N36_tdsp_state_1_),
		.A2(tdsp_state[0]),
		.B0(n_35),
		.B1(n_37),
		.Y(n_22));

	NAND3X1 i_41(
		.A(n_23),
		.B(n_72),
		.C(n_34),
		.Y(n_28));

	AOI21X1 i_5(
		.A0(bus_request),
		.A1(bus_grant),
		.B0(tdsp_state[0]),
		.Y(n_31));

	OAI21XL i_13(
		.A0(n_31),
		.A1(n_34),
		.B0(n_49),
		.Y(n_33));

	NAND2X1 i_2(
		.A(SPCASCAN_N31_tdsp_state_2_),
		.B(SPCASCAN_N36_tdsp_state_1_),
		.Y(n_34));

	NOR2BX1 i_1(
		.AN(SPCASCAN_N36_tdsp_state_1_),
		.B(SPCASCAN_N31_tdsp_state_2_),
		.Y(n_35));

	NOR2BX1 i_08999(
		.AN(bus_request),
		.B(bus_grant),
		.Y(n_36));

	NOR2X1 i_9(
		.A(n_36),
		.B(tdsp_state[0]),
		.Y(n_37));

	NOR2X1 i_4(
		.A(SPCASCAN_N36_tdsp_state_1_),
		.B(tdsp_state[0]),
		.Y(n_40));

	NAND4BXL i_17(
		.AN(n_57),
		.B(n_117),
		.C(n_102),
		.D(n_42),
		.Y(n_45));

	AOI22X1 i_24(
		.A0(n_35),
		.A1(n_36),
		.B0(SPCASCAN_N31_tdsp_state_2_),
		.B1(n_2818),
		.Y(n_47));

	NOR2X1 i_35(
		.A(n_36),
		.B(SPCASCAN_N31_tdsp_state_2_),
		.Y(n_48));

	SDFFRHQX1 tdsp_state_reg_0(
		.SI(BG_scan_in),
		.SE(scan_en),
		.D(n_33),
		.CK(clk),
		.RN(n_2820),
		.Q(tdsp_state[0]));

	SDFFRHQX1 tdsp_state_reg_1(
		.SI(FE_PT4_),
		.SE(scan_en),
		.D(n_28),
		.CK(clk),
		.RN(n_2820),
		.Q(SPCASCAN_N36_tdsp_state_1_));

	SDFFRHQX1 tdsp_state_reg_2(
		.SI(SPCASCAN_N32_two_cycle),
		.SE(scan_en),
		.D(n_27),
		.CK(clk),
		.RN(n_2820),
		.Q(SPCASCAN_N31_tdsp_state_2_));

	SDFFHQX1 samp_bio_reg(
		.SI(FE_PT1_),
		.SE(scan_en),
		.D(bio),
		.CK(clk),
		.Q(samp_bio));

	SDFFHQX1 samp_int_reg(
		.SI(phi_2),
		.SE(scan_en),
		.D(int),
		.CK(clk),
		.Q(SPCASCAN_N33_samp_int));

	SDFFRHQX1 phi_5_reg(
		.SI(tdsp_state[0]),
		.SE(scan_en),
		.D(n_2782),
		.CK(clk),
		.RN(n_2820),
		.Q(phi_5));

	OAI21XL i_598(
		.A0(n_24),
		.A1(n_2822),
		.B0(n_2784),
		.Y(n_2782));

	NAND3X1 i_599(
		.A(SPCASCAN_N31_tdsp_state_2_),
		.B(n_40),
		.C(n_24),
		.Y(n_2784));

	AOI21X1 i_37(
		.A0(n_48),
		.A1(n_2818),
		.B0(n_40),
		.Y(n_49));

	SDFFRHQX1 phi_4_reg(
		.SI(SPCASCAN_N34_two_cycle),
		.SE(scan_en),
		.D(n_2788),
		.CK(clk),
		.RN(n_2820),
		.Q(phi_4));

	OAI21XL i_605(
		.A0(n_24),
		.A1(n_2821),
		.B0(n_2790),
		.Y(n_2788));

	NAND3X1 i_606(
		.A(tdsp_state[0]),
		.B(n_35),
		.C(n_24),
		.Y(n_2790));

	NOR3X1 i_20(
		.A(SPCASCAN_N36_tdsp_state_1_),
		.B(SPCASCAN_N31_tdsp_state_2_),
		.C(tdsp_state[0]),
		.Y(n_57));

	SDFFRHQX1 phi_3_reg(
		.SI(FE_PT3_),
		.SE(scan_en),
		.D(n_2794),
		.CK(clk),
		.RN(n_2820),
		.Q(phi_3));

	OAI21XL i_612(
		.A0(n_22),
		.A1(n_2819),
		.B0(n_2797),
		.Y(n_2794));

	NAND2X1 i_614(
		.A(phi_3),
		.B(n_2819),
		.Y(n_2797));

	OR3XL i_23(
		.A(SPCASCAN_N31_tdsp_state_2_),
		.B(SPCASCAN_N36_tdsp_state_1_),
		.C(n_2818),
		.Y(n_72));

	SDFFRHQX1 phi_2_reg(
		.SI(phi_4),
		.SE(scan_en),
		.D(n_2800),
		.CK(clk),
		.RN(n_2820),
		.Q(phi_2));

	OAI21XL i_619(
		.A0(n_72),
		.A1(n_2819),
		.B0(n_2803),
		.Y(n_2800));

	NAND2X1 i_621(
		.A(phi_2),
		.B(n_2819),
		.Y(n_2803));

	NAND2X1 i_31(
		.A(n_35),
		.B(tdsp_state[0]),
		.Y(n_102));

	SDFFRHQX1 phi_1_reg(
		.SI(FE_PT2_),
		.SE(scan_en),
		.D(n_2806),
		.CK(clk),
		.RN(n_2820),
		.Q(phi_1));

	MX2X1 i_626(
		.S0(n_2819),
		.B(phi_1),
		.A(n_57),
		.Y(n_2806));

	NAND2X1 i_34(
		.A(SPCASCAN_N31_tdsp_state_2_),
		.B(n_40),
		.Y(n_117));

	SDFFRHQX1 phi_6_reg(
		.SI(SPCASCAN_N35_three_cycle),
		.SE(scan_en),
		.D(n_2812),
		.CK(clk),
		.RN(n_2820),
		.Q(BG_scan_out));

	OAI21XL i_633(
		.A0(n_42),
		.A1(n_2819),
		.B0(n_2815),
		.Y(n_2812));

	NAND2X1 i_635(
		.A(phi_6),
		.B(n_2819),
		.Y(n_2815));

	NAND3BX1 i_36(
		.AN(SPCASCAN_N36_tdsp_state_1_),
		.B(SPCASCAN_N31_tdsp_state_2_),
		.C(tdsp_state[0]),
		.Y(n_42));

	INVX1 i_682(
		.A(tdsp_state[0]),
		.Y(n_2818));

	INVX1 i_683(
		.A(n_24),
		.Y(n_2819));

	INVX1 i_684(
		.A(reset),
		.Y(n_2820));

	INVX1 i_685(
		.A(phi_4),
		.Y(n_2821));

	INVX1 i_686(
		.A(phi_5),
		.Y(n_2822));

endmodule
module tdsp_core(
		clk,
		reset,
		as,
		read,
		write,
		address,
		t_data_in,
		t_data_out,
		p_read,
		p_address,
		rom_data_in,
		bus_grant,
		bus_request,
		port_as,
		port_address,
		port_pad_data_in,
		port_pad_data_out,
		bio,
		int,
		scan_en,
		BG_scan_in,
		BG_scan_out,
	SPCASCAN_N1_p_data_out_13_,
	SPCASCAN_N2_low_mag_8_,
	SPCASCAN_N3_port_data_out_0_,
	SPCASCAN_N4_low_mag_3_,
	SPCASCAN_N5_port_data_out_1_,
	FE_PT1_,
	SPCASCAN_N22_data_out_0_,
	SPCASCAN_N24_t_sel_7,
	SPCASCAN_N25_data_out_12_,
	SPCASCAN_N26_spi_sr_0_,
	SPCASCAN_N27_port_data_out_11_,
	n_7862);
   output SPCASCAN_N1_p_data_out_13_;
   input SPCASCAN_N2_low_mag_8_;
   output SPCASCAN_N3_port_data_out_0_;
   input SPCASCAN_N4_low_mag_3_;
   output SPCASCAN_N5_port_data_out_1_;
   input FE_PT1_;
   output SPCASCAN_N22_data_out_0_;
   input SPCASCAN_N24_t_sel_7;
   output SPCASCAN_N25_data_out_12_;
   input SPCASCAN_N26_spi_sr_0_;
   output SPCASCAN_N27_port_data_out_11_;
   input n_7862;

	input clk;
	input reset;
	output as;
	output read;
	output write;
	output [7:0] address;
	input [15:0] t_data_in;
	output [15:0] t_data_out;
	output p_read;
	output [8:0] p_address;
	input [15:0] rom_data_in;
	input bus_grant;
	output bus_request;
	output port_as;
	output [2:0] port_address;
	input [15:0] port_pad_data_in;
	output [15:0] port_pad_data_out;
	input bio;
	input int;
	input scan_en;
	input BG_scan_in;
	output BG_scan_out;

	wire [15:0] data_out;
	wire [15:0] data_in;
	wire [15:0] ir;
	wire [15:0] port_data_in;
	wire [2:0] port_addrs_in;
	wire [8:0] p_addrs_in;
	wire [2:0] sel_op_b;
	wire [2:0] sel_op_a;
	wire [15:0] top;
	wire [31:0] p;
	wire [15:0] ar1;
	wire [15:0] ar0;
	wire [15:0] port_data_out;
	wire [15:0] p_data_out;
	wire [7:0] addrs_in;
	wire [15:0] decode;
	wire [15:0] ar;
	wire [15:0] mdr;
	wire [31:0] mpy_result;
	wire [32:0] alu_result;
	wire [3:0] alu_cmd;
	wire [31:0] opb;
	wire [31:0] opa;



	BUFX1 i_10181(
		.A(opa[11]),
		.Y(n_7285));

	BUFX2 i_10177(
		.A(opa[8]),
		.Y(n_7280));

	BUFX2 i_10173(
		.A(opa[9]),
		.Y(n_7275));

	BUFX1 i_10155(
		.A(opa[12]),
		.Y(n_7252));

	CLKBUFX2 i_10149(
		.A(opa[13]),
		.Y(n_7244));

	BUFX1 i_10084(
		.A(ir[14]),
		.Y(n_7149));

	CLKBUFX3 i_9488(
		.A(\nbus_642[1] ),
		.Y(address[1]));

	CLKBUFX3 i_9479(
		.A(ir[8]),
		.Y(n_6217));

	tdsp_core_mach TDSP_CORE_MACH_INST(
		.samp_bio(samp_bio),
		.phi_1(phi_1),
		.phi_3(phi_3),
		.phi_4(phi_4),
		.phi_5(phi_5),
		.phi_6(phi_6),
		.reset(reset),
		.clk(clk),
		.bus_request(bus_request),
		.bus_grant(bus_grant),
		.bio(bio),
		.int(int),
		.scan_en(scan_en),
		.BG_scan_in(dec_read_data),
		.BG_scan_out(n_7866),
	.FE_PT1_(data_out[11]),
	.SPCASCAN_N31_tdsp_state_2_(SPCASCAN_N31_tdsp_state_2_),
	.SPCASCAN_N32_two_cycle(SPCASCAN_N32_two_cycle),
	.FE_PT2_(\acc[21] ),
	.SPCASCAN_N33_samp_int(SPCASCAN_N33_samp_int),
	.SPCASCAN_N34_two_cycle(SPCASCAN_N34_two_cycle),
	.SPCASCAN_N35_three_cycle(SPCASCAN_N35_three_cycle),
	.FE_PT3_(\acc[19] ),
	.SPCASCAN_N36_tdsp_state_1_(SPCASCAN_N36_tdsp_state_1_),
	.FE_PT4_(\acc[20] ));

	prog_bus_mach PROG_BUS_MACH_INST(
		.clk(clk),
		.reset(reset),
		.read(p_read),
		.address(p_address),
		.data_out({ p_data_out[15], p_data_out[14], SPCASCAN_N1_p_data_out_13_,
	p_data_out[12], p_data_out[11], p_data_out[10],
	p_data_out[9], p_data_out[8], p_data_out[7],
	p_data_out[6], p_data_out[5], p_data_out[4],
	p_data_out[3], p_data_out[2], p_data_out[1],
	p_data_out[0]}),
		.pad_data_in(rom_data_in),
		.addrs_in(p_addrs_in),
		.read_cycle(read_prog),
		.go(go_prog),
		.scan_en(scan_en),
		.BG_scan_in(n_7866),
		.BG_scan_out(n_7867),
	.FE_PT1_(port_data_out[5]),
	.FE_PT2_(p[24]),
	.SPCASCAN_N6_present_state_2_(SPCASCAN_N6_present_state_2_),
	.FE_PT3_(p[29]),
	.SPCASCAN_N7_present_state_1_(SPCASCAN_N7_present_state_1_),
	.FE_PT4_(data_out[4]),
	.FE_PT5_(\pc[1] ));

	port_bus_mach PORT_BUS_MACH_INST(
		.clk(clk),
		.reset(reset),
		.address(port_address),
		.data_in(port_data_in),
		.data_out({ port_data_out[15], port_data_out[14], port_data_out[13],
	port_data_out[12], SPCASCAN_N27_port_data_out_11_, port_data_out[10],
	port_data_out[9], port_data_out[8], port_data_out[7],
	port_data_out[6], port_data_out[5], port_data_out[4],
	port_data_out[3], port_data_out[2], SPCASCAN_N5_port_data_out_1_,
	SPCASCAN_N3_port_data_out_0_}),
		.pad_data_in(port_pad_data_in),
		.pad_data_out(port_pad_data_out),
		.addrs_in(port_addrs_in),
		.read_cycle(read_port),
		.go(go_port),
		.as(port_as),
		.scan_en(scan_en),
		.BG_scan_in(n_7867),
		.BG_scan_out(n_7868),
	.SPCASCAN_N2_low_mag_8_(SPCASCAN_N2_low_mag_8_),
	.SPCASCAN_N4_low_mag_3_(SPCASCAN_N4_low_mag_3_),
	.p_read(p_read),
	.SPCASCAN_N26_spi_sr_0_(SPCASCAN_N26_spi_sr_0_),
	.FE_PT1_(data_out[10]),
	.SPCASCAN_N28_read(SPCASCAN_N28_read),
	.FE_PT2_(ar0[0]),
	.FE_PT3_(ar0[13]),
	.SPCASCAN_N29_present_state_1_(SPCASCAN_N29_present_state_1_),
	.FE_PT4_(ar0[3]),
	.FE_PT5_(ar1[0]),
	.SPCASCAN_N30_ov(SPCASCAN_N30_ov));

	alu_32 ALU_32_INST(
		.ovm(ovm),
		.op_a({
		opa[31],
		opa[30],
		opa[29],
		opa[28],
		opa[27],
		opa[26],
		opa[25],
		opa[24],
		opa[23],
		opa[22],
		opa[21],
		opa[20],
		opa[19],
		opa[18],
		opa[17],
		opa[16],
		opa[15],
		opa[14],
		n_7244,
		n_7252,
		n_7285,
		opa[10],
		n_7275,
		n_7280,
		opa[7],
		opa[6],
		opa[5],
		opa[4],
		opa[3],
		opa[2],
		opa[1],
		opa[0]}),
		.op_b(opb),
		.result(alu_result),
		.cmd(alu_cmd));

	mult_32 MPY_32_INST(
		.op_a({
		opa[15],
		opa[14],
		opa[13],
		opa[12],
		opa[11],
		opa[10],
		opa[9],
		opa[8],
		opa[7],
		opa[6],
		opa[5],
		opa[4],
		opa[3],
		opa[2],
		opa[1],
		opa[0]}),
		.op_b({
		opb[15],
		opb[14],
		opb[13],
		opb[12],
		opb[11],
		opb[10],
		opb[9],
		opb[8],
		opb[7],
		opb[6],
		opb[5],
		opb[4],
		opb[3],
		opb[2],
		opb[1],
		opb[0]}),
		.result(mpy_result));

	accum_stat ACCUM_STAT_INST(
		.accum({
		UNCONNECTED_000,
		\acc[31] ,
		\acc[30] ,
		\acc[29] ,
		\acc[28] ,
		\acc[27] ,
		\acc[26] ,
		\acc[25] ,
		\acc[24] ,
		\acc[23] ,
		\acc[22] ,
		\acc[21] ,
		\acc[20] ,
		\acc[19] ,
		\acc[18] ,
		\acc[17] ,
		\acc[16] ,
		\acc[15] ,
		\acc[14] ,
		\acc[13] ,
		\acc[12] ,
		\acc[11] ,
		\acc[10] ,
		\acc[9] ,
		\acc[8] ,
		\acc[7] ,
		\acc[6] ,
		\acc[5] ,
		\acc[4] ,
		\acc[3] ,
		\acc[2] ,
		\acc[1] ,
		\acc[0] }),
		.ar(ar),
		.bio(samp_bio),
		.gez(gez),
		.gz(gz),
		.nz(nz),
		.lz(lz),
		.lez(lez),
		.arnz(arnz),
		.bioz(bioz));

	execute_i EXECUTE_INST(
		.clk(clk),
		.reset(reset),
		.phi_1(phi_1),
		.phi_3(phi_3),
		.phi_4(phi_4),
		.phi_5(phi_5),
		.phi_6(phi_6),
		.gez(gez),
		.gz(gz),
		.nz(nz),
		.lz(lz),
		.lez(lez),
		.arnz(arnz),
		.bioz(bioz),
		.alu_result(alu_result),
		.mpy_result(mpy_result),
		.mdr(mdr),
		.ir({
		ir[15],
		n_7149,
		ir[13],
		ir[12],
		ir[11],
		ir[10],
		ir[9],
		n_6217,
		ir[7],
		ir[6],
		ir[5],
		ir[4],
		ir[3],
		ir[2],
		ir[1],
		ir[0]}),
		.decode(decode),
		.ar(ar),
		.skip_one(skip_one),
		.pc_acc(pc_acc),
		.dmov_inc(dmov_inc),
		.dp(dp),
		.arp(arp),
		.ar0(ar0),
		.ar1(ar1),
		.pc({
		UNCONNECTED_001,
		UNCONNECTED_002,
		UNCONNECTED_003,
		UNCONNECTED_004,
		UNCONNECTED_005,
		UNCONNECTED_006,
		UNCONNECTED_007,
		\pc[8] ,
		\pc[7] ,
		\pc[6] ,
		\pc[5] ,
		\pc[4] ,
		\pc[3] ,
		\pc[2] ,
		\pc[1] ,
		\pc[0] }),
		.acc({
		UNCONNECTED_008,
		\acc[31] ,
		\acc[30] ,
		\acc[29] ,
		\acc[28] ,
		\acc[27] ,
		\acc[26] ,
		\acc[25] ,
		\acc[24] ,
		\acc[23] ,
		\acc[22] ,
		\acc[21] ,
		\acc[20] ,
		\acc[19] ,
		\acc[18] ,
		\acc[17] ,
		\acc[16] ,
		\acc[15] ,
		\acc[14] ,
		\acc[13] ,
		\acc[12] ,
		\acc[11] ,
		\acc[10] ,
		\acc[9] ,
		\acc[8] ,
		\acc[7] ,
		\acc[6] ,
		\acc[5] ,
		\acc[4] ,
		\acc[3] ,
		\acc[2] ,
		\acc[1] ,
		\acc[0] }),
		.p(p),
		.top(top),
		.alu_cmd(alu_cmd),
		.sel_op_a(sel_op_a),
		.sel_op_b(sel_op_b),
		.read_prog(enc_read_prog),
		.go_prog(enc_go_prog),
		.read_data(enc_read_data),
		.go_data(enc_go_data),
		.read_port(enc_read_port),
		.go_port(enc_go_port),
		.ovm(ovm),
		.scan_en(scan_en),
		.BG_scan_in(n_7868),
		.BG_scan_out(n_7869),
	.SPCASCAN_N6_present_state_2_(SPCASCAN_N6_present_state_2_),
	.SPCASCAN_N7_present_state_1_(SPCASCAN_N7_present_state_1_),
	.FE_PT1_(data_out[1]),
	.SPCASCAN_N23_done(SPCASCAN_N23_done),
	.SPCASCAN_N28_read(SPCASCAN_N28_read),
	.port_as(port_as),
	.FE_PT2_(ir[8]),
	.dec_go_port(dec_go_port),
	.SPCASCAN_N29_present_state_1_(SPCASCAN_N29_present_state_1_),
	.FE_PT3_(port_data_out[13]),
	.FE_PT4_(port_data_out[14]),
	.SPCASCAN_N30_ov(SPCASCAN_N30_ov),
	.SPCASCAN_N31_tdsp_state_2_(SPCASCAN_N31_tdsp_state_2_),
	.SPCASCAN_N32_two_cycle(SPCASCAN_N32_two_cycle),
	.SPCASCAN_N33_samp_int(SPCASCAN_N33_samp_int),
	.n_7866(n_7866),
	.SPCASCAN_N35_three_cycle(SPCASCAN_N35_three_cycle),
	.dec_go_data(dec_go_data),
	.dec_go_prog(dec_go_prog),
	.SPCASCAN_N36_tdsp_state_1_(SPCASCAN_N36_tdsp_state_1_),
	.n_7862(n_7862));

	decode_i DECODE_INST(
		.clk(clk),
		.reset(reset),
		.phi_3(phi_3),
		.phi_6(phi_6),
		.decode(decode),
		.p_data_out({ p_data_out[15], p_data_out[14], SPCASCAN_N1_p_data_out_13_,
	p_data_out[12], p_data_out[11], p_data_out[10],
	p_data_out[9], p_data_out[8], p_data_out[7],
	p_data_out[6], p_data_out[5], p_data_out[4],
	p_data_out[3], p_data_out[2], p_data_out[1],
	p_data_out[0]}),
		.ir(ir),
		.skip_one(skip_one),
		.read_prog(dec_read_prog),
		.go_prog(dec_go_prog),
		.read_data(dec_read_data),
		.go_data(dec_go_data),
		.read_port(dec_read_port),
		.go_port(dec_go_port),
		.scan_en(scan_en),
		.BG_scan_in(n_7869),
		.BG_scan_out(n_7870),
	.FE_PT1_(ar0[15]),
	.FE_PT2_(ar1[11]),
	.FE_PT3_(\pc[8] ),
	.FE_PT4_(\pc[4] ),
	.FE_PT5_(\pc[3] ),
	.FE_PT6_(\pc[7] ),
	.FE_PT7_(top[11]),
	.FE_PT8_(top[3]),
	.arp(arp),
	.pc_acc(pc_acc),
	.SPCASCAN_N34_two_cycle(SPCASCAN_N34_two_cycle),
	.enc_read_port(enc_read_port),
	.UNCONNECTED_006(UNCONNECTED_006),
	.enc_go_data(enc_go_data),
	.enc_read_data(enc_read_data));

	tdsp_core_glue TDSP_CORE_GLUE_INST(
		.addrs_in(addrs_in),
		.data_in(data_in),
		.p_addrs_in(p_addrs_in),
		.port_addrs_in(port_addrs_in),
		.port_data_in(port_data_in),
		.ar(ar),
		.go_prog(go_prog),
		.read_prog(read_prog),
		.go_data(go_data),
		.read_data(read_data),
		.go_port(go_port),
		.read_port(read_port),
		.pc_acc(pc_acc),
		.arp(arp),
		.ar1(ar1),
		.ar0(ar0),
		.dp(dp),
		.ir({
		ir[15],
		ir[14],
		ir[13],
		ir[12],
		ir[11],
		ir[10],
		ir[9],
		n_6217,
		ir[7],
		ir[6],
		ir[5],
		ir[4],
		ir[3],
		ir[2],
		ir[1],
		ir[0]}),
		.opa(opa),
		.opb(opb),
		.mdr(mdr),
		.acc({
		UNCONNECTED_009,
		\acc[31] ,
		\acc[30] ,
		\acc[29] ,
		\acc[28] ,
		\acc[27] ,
		\acc[26] ,
		\acc[25] ,
		\acc[24] ,
		\acc[23] ,
		\acc[22] ,
		\acc[21] ,
		\acc[20] ,
		\acc[19] ,
		\acc[18] ,
		\acc[17] ,
		\acc[16] ,
		\acc[15] ,
		\acc[14] ,
		\acc[13] ,
		\acc[12] ,
		\acc[11] ,
		\acc[10] ,
		\acc[9] ,
		\acc[8] ,
		\acc[7] ,
		\acc[6] ,
		\acc[5] ,
		\acc[4] ,
		\acc[3] ,
		\acc[2] ,
		\acc[1] ,
		\acc[0] }),
		.pc({
		UNCONNECTED_010,
		UNCONNECTED_011,
		UNCONNECTED_012,
		UNCONNECTED_013,
		UNCONNECTED_014,
		UNCONNECTED_015,
		UNCONNECTED_016,
		\pc[8] ,
		\pc[7] ,
		\pc[6] ,
		\pc[5] ,
		\pc[4] ,
		\pc[3] ,
		\pc[2] ,
		\pc[1] ,
		\pc[0] }),
		.data_out({ data_out[15], data_out[14], data_out[13],
	SPCASCAN_N25_data_out_12_, data_out[11], data_out[10],
	data_out[9], data_out[8], data_out[7],
	data_out[6], data_out[5], data_out[4],
	data_out[3], data_out[2], data_out[1],
	SPCASCAN_N22_data_out_0_}),
		.p_data_out({ p_data_out[15], p_data_out[14], SPCASCAN_N1_p_data_out_13_,
	p_data_out[12], p_data_out[11], p_data_out[10],
	p_data_out[9], p_data_out[8], p_data_out[7],
	p_data_out[6], p_data_out[5], p_data_out[4],
	p_data_out[3], p_data_out[2], p_data_out[1],
	p_data_out[0]}),
		.port_data_out({ port_data_out[15], port_data_out[14], port_data_out[13],
	port_data_out[12], SPCASCAN_N27_port_data_out_11_, port_data_out[10],
	port_data_out[9], port_data_out[8], port_data_out[7],
	port_data_out[6], port_data_out[5], port_data_out[4],
	port_data_out[3], port_data_out[2], SPCASCAN_N5_port_data_out_1_,
	SPCASCAN_N3_port_data_out_0_}),
		.top(top),
		.p(p),
		.sel_op_a(sel_op_a),
		.sel_op_b(sel_op_b),
		.dec_go_prog(dec_go_prog),
		.enc_go_prog(enc_go_prog),
		.dec_read_prog(dec_read_prog),
		.enc_read_prog(enc_read_prog),
		.dec_go_data(dec_go_data),
		.enc_go_data(enc_go_data),
		.dec_read_data(dec_read_data),
		.enc_read_data(enc_read_data),
		.dec_go_port(dec_go_port),
		.enc_go_port(enc_go_port),
		.dec_read_port(dec_read_port),
		.enc_read_port(enc_read_port),
		.dmov_inc(dmov_inc));

	data_bus_mach DATA_BUS_MACH_INST(
		.clk(clk),
		.reset(reset),
		.read(read),
		.write(write),
		.address({
		address[7],
		address[6],
		address[5],
		address[4],
		address[3],
		address[2],
		\nbus_642[1] ,
		address[0]}),
		.data_in(data_in),
		.data_out({ data_out[15], data_out[14], data_out[13],
	SPCASCAN_N25_data_out_12_, data_out[11], data_out[10],
	data_out[9], data_out[8], data_out[7],
	data_out[6], data_out[5], data_out[4],
	data_out[3], data_out[2], data_out[1],
	SPCASCAN_N22_data_out_0_}),
		.pad_data_in(t_data_in),
		.pad_data_out(t_data_out),
		.addrs_in(addrs_in),
		.read_cycle(read_data),
		.go(go_data),
		.as(as),
		.bus_request(bus_request),
		.bus_grant(bus_grant),
		.scan_en(scan_en),
		.BG_scan_in(read),
		.BG_scan_out(BG_scan_out),
	.FE_PT1_(FE_PT1_),
	.n_7867(n_7867),
	.FE_PT2_(\pc[0] ),
	.SPCASCAN_N23_done(SPCASCAN_N23_done),
	.SPCASCAN_N24_t_sel_7(SPCASCAN_N24_t_sel_7),
	.FE_PT3_(port_data_out[7]),
	.samp_bio(samp_bio),
	.FE_PT4_(ar1[9]));

endmodule
module ADDFHX1 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule
module ADDFHX2 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule
module ADDFHX4 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule
module ADDFHXL ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule
module ADDFX1 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule
module ADDFX2 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule
module ADDFX4 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule
module ADDFXL ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule
module ADDHX1 ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule
module ADDHX2 ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule
module ADDHX4 ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule
module ADDHXL ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule
module AFCSHCINX2 ( CS, A, B, CI0N, CI1N, S, CO0, CO1);
    input		CS ;
    input		A ;
    input		B ;
    input		CI0N ;
    input		CI1N ;
    output		S ;
    output		CO0 ;
    output		CO1 ;

endmodule
module AFCSHCINX4 ( CS, A, B, CI0N, CI1N, S, CO0, CO1);
    input		CS ;
    input		A ;
    input		B ;
    input		CI0N ;
    input		CI1N ;
    output		S ;
    output		CO0 ;
    output		CO1 ;

endmodule
module AFCSHCONX2 ( CS, A, B, CI0, CI1, S, CO0N, CO1N);
    input		CS ;
    input		A ;
    input		B ;
    input		CI0 ;
    input		CI1 ;
    output		S ;
    output		CO0N ;
    output		CO1N ;

endmodule
module AFCSHCONX4 ( CS, A, B, CI0, CI1, S, CO0N, CO1N);
    input		CS ;
    input		A ;
    input		B ;
    input		CI0 ;
    input		CI1 ;
    output		S ;
    output		CO0N ;
    output		CO1N ;

endmodule
module AFHCINX2 ( A, B, CIN, S, CO);
    input		A ;
    input		B ;
    input		CIN ;
    output		S ;
    output		CO ;

endmodule
module AFHCINX4 ( A, B, CIN, S, CO);
    input		A ;
    input		B ;
    input		CIN ;
    output		S ;
    output		CO ;

endmodule
module AFHCONX2 ( A, B, CI, S, CON);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CON ;

endmodule
module AFHCONX4 ( A, B, CI, S, CON);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CON ;

endmodule
module AHHCINX2 ( A, CIN, S, CO);
    input		A ;
    input		CIN ;
    output		S ;
    output		CO ;

endmodule
module AHHCINX4 ( A, CIN, S, CO);
    input		A ;
    input		CIN ;
    output		S ;
    output		CO ;

endmodule
module AHHCONX2 ( A, CI, S, CON);
    input		A ;
    input		CI ;
    output		S ;
    output		CON ;

endmodule
module AHHCONX4 ( A, CI, S, CON);
    input		A ;
    input		CI ;
    output		S ;
    output		CON ;

endmodule
module AND2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module AND2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module AND2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module AND2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module AND3X1 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module AND3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module AND3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module AND3XL ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module AND4X1 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module AND4X2 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module AND4X4 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module AND4XL ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module AOI211X1 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule
module AOI211X2 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule
module AOI211X4 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule
module AOI211XL ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule
module AOI21X1 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule
module AOI21X2 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule
module AOI21X4 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule
module AOI21XL ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule
module AOI221X1 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule
module AOI221X2 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule
module AOI221X4 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule
module AOI221XL ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule
module AOI222X1 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule
module AOI222X2 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule
module AOI222X4 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule
module AOI222XL ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule
module AOI22X1 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI22X2 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI22X4 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI22XL ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI2BB1X1 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule
module AOI2BB1X2 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule
module AOI2BB1X4 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule
module AOI2BB1XL ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule
module AOI2BB2X1 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI2BB2X2 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI2BB2X4 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI2BB2XL ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI31X1 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule
module AOI31X2 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule
module AOI31X4 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule
module AOI31XL ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule
module AOI32X1 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI32X2 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI32X4 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI32XL ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module AOI33X1 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule
module AOI33X2 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule
module AOI33X4 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule
module AOI33XL ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule
module BENCX1 ( M2, M1, M0, A, S, X2);
    input		M2 ;
    input		M1 ;
    input		M0 ;
    output		A ;
    output		S ;
    output		X2 ;

endmodule
module BENCX2 ( M2, M1, M0, A, S, X2);
    input		M2 ;
    input		M1 ;
    input		M0 ;
    output		A ;
    output		S ;
    output		X2 ;

endmodule
module BENCX4 ( M2, M1, M0, A, S, X2);
    input		M2 ;
    input		M1 ;
    input		M0 ;
    output		A ;
    output		S ;
    output		X2 ;

endmodule
module BMXX1 ( X2, M0, A, S, M1, PP);
    input		X2 ;
    input		M0 ;
    input		A ;
    input		S ;
    input		M1 ;
    output		PP ;

endmodule
module BUFX1 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module BUFX12 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module BUFX16 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module BUFX2 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module BUFX20 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module BUFX3 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module BUFX4 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module BUFX8 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module BUFXL ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFX1 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFX12 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFX16 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFX2 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFX20 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFX3 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFX4 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFX8 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKBUFXL ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVX1 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVX12 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVX16 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVX2 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVX20 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVX3 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVX4 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVX8 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CLKINVXL ( A, Y);
    input		A ;
    output		Y ;

endmodule
module CMPR22X1 ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule
module CMPR32X1 ( A, B, C, S, CO);
    input		A ;
    input		B ;
    input		C ;
    output		S ;
    output		CO ;

endmodule
module CMPR42X1 ( A, B, C, D, ICI, S, ICO, CO);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    input		ICI ;
    output		S ;
    output		ICO ;
    output		CO ;

endmodule
module CMPR42X2 ( A, B, C, D, ICI, S, ICO, CO);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    input		ICI ;
    output		S ;
    output		ICO ;
    output		CO ;

endmodule
module DFFHQX1 ( D, CK, Q);
    input		D ;
    input		CK ;
    output		Q ;

endmodule
module DFFHQX2 ( D, CK, Q);
    input		D ;
    input		CK ;
    output		Q ;

endmodule
module DFFHQX4 ( D, CK, Q);
    input		D ;
    input		CK ;
    output		Q ;

endmodule
module DFFHQXL ( D, CK, Q);
    input		D ;
    input		CK ;
    output		Q ;

endmodule
module DFFNRX1 ( D, CKN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNRX2 ( D, CKN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNRX4 ( D, CKN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNRXL ( D, CKN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNSRX1 ( D, CKN, SN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNSRX2 ( D, CKN, SN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNSRX4 ( D, CKN, SN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNSRXL ( D, CKN, SN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNSX1 ( D, CKN, SN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNSX2 ( D, CKN, SN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNSX4 ( D, CKN, SN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNSXL ( D, CKN, SN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNX1 ( D, CKN, Q, QN);
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNX2 ( D, CKN, Q, QN);
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNX4 ( D, CKN, Q, QN);
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule
module DFFNXL ( D, CKN, Q, QN);
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule
module DFFRHQX1 ( D, CK, RN, Q);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule
module DFFRHQX2 ( D, CK, RN, Q);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule
module DFFRHQX4 ( D, CK, RN, Q);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule
module DFFRHQXL ( D, CK, RN, Q);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule
module DFFRX1 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFRX2 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFRX4 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFRXL ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFSHQX1 ( D, CK, SN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule
module DFFSHQX2 ( D, CK, SN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule
module DFFSHQX4 ( D, CK, SN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule
module DFFSHQXL ( D, CK, SN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule
module DFFSRHQX1 ( D, CK, SN, RN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule
module DFFSRHQX2 ( D, CK, SN, RN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule
module DFFSRHQX4 ( D, CK, SN, RN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule
module DFFSRHQXL ( D, CK, SN, RN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule
module DFFSRX1 ( D, CK, SN, RN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFSRX2 ( D, CK, SN, RN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFSRX4 ( D, CK, SN, RN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFSRXL ( D, CK, SN, RN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFSX1 ( D, CK, SN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module DFFSX2 ( D, CK, SN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module DFFSX4 ( D, CK, SN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module DFFSXL ( D, CK, SN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module DFFTRX1 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFTRX2 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFTRX4 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFTRXL ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module DFFX1 ( D, CK, Q, QN);
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module DFFX2 ( D, CK, Q, QN);
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module DFFX4 ( D, CK, Q, QN);
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module DFFXL ( D, CK, Q, QN);
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module DLY1X1 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module DLY2X1 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module DLY3X1 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module DLY4X1 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module EDFFTRX1 ( D, CK, E, RN, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module EDFFTRX2 ( D, CK, E, RN, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module EDFFTRX4 ( D, CK, E, RN, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module EDFFTRXL ( D, CK, E, RN, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module EDFFX1 ( D, CK, E, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule
module EDFFX2 ( D, CK, E, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule
module EDFFX4 ( D, CK, E, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule
module EDFFXL ( D, CK, E, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule
module HOLDX1 ( Y);
    inout		Y ;

endmodule
module INVX1 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module INVX12 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module INVX16 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module INVX2 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module INVX20 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module INVX3 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module INVX4 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module INVX8 ( A, Y);
    input		A ;
    output		Y ;

endmodule
module INVXL ( A, Y);
    input		A ;
    output		Y ;

endmodule
module JKFFRX1 ( J, K, CK, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFRX2 ( J, K, CK, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFRX4 ( J, K, CK, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFRXL ( J, K, CK, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFSRX1 ( J, K, CK, SN, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFSRX2 ( J, K, CK, SN, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFSRX4 ( J, K, CK, SN, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFSRXL ( J, K, CK, SN, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFSX1 ( J, K, CK, SN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFSX2 ( J, K, CK, SN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFSX4 ( J, K, CK, SN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFSXL ( J, K, CK, SN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module JKFFX1 ( J, K, CK, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module JKFFX2 ( J, K, CK, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module JKFFX4 ( J, K, CK, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module JKFFXL ( J, K, CK, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module MX2X1 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MX2X2 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MX2X4 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MX2XL ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MX4X1 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MX4X2 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MX4X4 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MX4XL ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MXI2X1 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MXI2X2 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MXI2X4 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MXI2XL ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MXI4X1 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MXI4X2 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MXI4X4 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module MXI4XL ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule
module NAND2BX1 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule
module NAND2BX2 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule
module NAND2BX4 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule
module NAND2BXL ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule
module NAND2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module NAND2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module NAND2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module NAND2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module NAND3BX1 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NAND3BX2 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NAND3BX4 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NAND3BXL ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NAND3X1 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NAND3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NAND3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NAND3XL ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NAND4BBX1 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4BBX2 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4BBX4 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4BBXL ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4BX1 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4BX2 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4BX4 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4BXL ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4X1 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4X2 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4X4 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NAND4XL ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR2BX1 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule
module NOR2BX2 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule
module NOR2BX4 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule
module NOR2BXL ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule
module NOR2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module NOR2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module NOR2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module NOR2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module NOR3BX1 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NOR3BX2 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NOR3BX4 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NOR3BXL ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NOR3X1 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NOR3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NOR3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NOR3XL ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module NOR4BBX1 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4BBX2 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4BBX4 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4BBXL ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4BX1 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4BX2 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4BX4 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4BXL ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4X1 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4X2 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4X4 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module NOR4XL ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module OAI211X1 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule
module OAI211X2 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule
module OAI211X4 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule
module OAI211XL ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule
module OAI21X1 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule
module OAI21X2 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule
module OAI21X4 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule
module OAI21XL ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule
module OAI221X1 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule
module OAI221X2 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule
module OAI221X4 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule
module OAI221XL ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule
module OAI222X1 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule
module OAI222X2 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule
module OAI222X4 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule
module OAI222XL ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule
module OAI22X1 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI22X2 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI22X4 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI22XL ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI2BB1X1 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule
module OAI2BB1X2 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule
module OAI2BB1X4 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule
module OAI2BB1XL ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule
module OAI2BB2X1 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI2BB2X2 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI2BB2X4 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI2BB2XL ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI31X1 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule
module OAI31X2 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule
module OAI31X4 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule
module OAI31XL ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule
module OAI32X1 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI32X2 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI32X4 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI32XL ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule
module OAI33X1 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule
module OAI33X2 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule
module OAI33X4 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule
module OAI33XL ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule
module OR2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module OR2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module OR2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module OR2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module OR3X1 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module OR3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module OR3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module OR3XL ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module OR4X1 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module OR4X2 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module OR4X4 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module OR4XL ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule
module RF1R1WX2 ( WW, WB, RW, RWN, RB);
    input		WW ;
    input		WB ;
    input		RW ;
    input		RWN ;
    output		RB ;

endmodule
module RF2R1WX2 ( WB, WW, R1W, R2W, R1B, R2B);
    input		WB ;
    input		WW ;
    input		R1W ;
    input		R2W ;
    output		R1B ;
    output		R2B ;

endmodule
module RFRDX1 ( RB, BRB);
    input		RB ;
    output		BRB ;

endmodule
module RFRDX2 ( RB, BRB);
    input		RB ;
    output		BRB ;

endmodule
module RFRDX4 ( RB, BRB);
    input		RB ;
    output		BRB ;

endmodule
module SDFFHQX1 ( SI, SE, D, CK, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;

endmodule
module SDFFHQX2 ( SI, SE, D, CK, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;

endmodule
module SDFFHQX4 ( SI, SE, D, CK, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;

endmodule
module SDFFHQXL ( SI, SE, D, CK, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;

endmodule
module SDFFNRX1 ( SI, SE, D, CKN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNRX2 ( SI, SE, D, CKN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNRX4 ( SI, SE, D, CKN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNRXL ( SI, SE, D, CKN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNSRX1 ( SI, SE, D, CKN, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNSRX2 ( SI, SE, D, CKN, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNSRX4 ( SI, SE, D, CKN, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNSRXL ( SI, SE, D, CKN, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNSX1 ( SI, SE, D, CKN, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNSX2 ( SI, SE, D, CKN, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNSX4 ( SI, SE, D, CKN, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNSXL ( SI, SE, D, CKN, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNX1 ( SI, SE, D, CKN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNX2 ( SI, SE, D, CKN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNX4 ( SI, SE, D, CKN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFNXL ( SI, SE, D, CKN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFRHQX1 ( SI, SE, D, CK, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule
module SDFFRHQX2 ( SI, SE, D, CK, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule
module SDFFRHQX4 ( SI, SE, D, CK, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule
module SDFFRHQXL ( SI, SE, D, CK, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule
module SDFFRX1 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFRX2 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFRX4 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFRXL ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFSHQX1 ( SI, SE, D, CK, SN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule
module SDFFSHQX2 ( SI, SE, D, CK, SN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule
module SDFFSHQX4 ( SI, SE, D, CK, SN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule
module SDFFSHQXL ( SI, SE, D, CK, SN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule
module SDFFSRHQX1 ( SI, SE, D, CK, SN, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule
module SDFFSRHQX2 ( SI, SE, D, CK, SN, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule
module SDFFSRHQX4 ( SI, SE, D, CK, SN, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule
module SDFFSRHQXL ( SI, SE, D, CK, SN, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule
module SDFFSRX1 ( SI, SE, D, CK, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFSRX2 ( SI, SE, D, CK, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFSRX4 ( SI, SE, D, CK, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFSRXL ( SI, SE, D, CK, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFSX1 ( SI, SE, D, CK, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFSX2 ( SI, SE, D, CK, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFSX4 ( SI, SE, D, CK, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFSXL ( SI, SE, D, CK, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFTRX1 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFTRX2 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFTRX4 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFTRXL ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SDFFX1 ( SI, SE, D, CK, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module SDFFX2 ( SI, SE, D, CK, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module SDFFX4 ( SI, SE, D, CK, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module SDFFXL ( SI, SE, D, CK, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule
module SEDFFHQX1 ( SI, SE, D, CK, E, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;

endmodule
module SEDFFHQX2 ( SI, SE, D, CK, E, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;

endmodule
module SEDFFHQX4 ( SI, SE, D, CK, E, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;

endmodule
module SEDFFHQXL ( SI, SE, D, CK, E, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;

endmodule
module SEDFFTRX1 ( SI, SE, D, CK, E, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SEDFFTRX2 ( SI, SE, D, CK, E, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SEDFFTRX4 ( SI, SE, D, CK, E, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SEDFFTRXL ( SI, SE, D, CK, E, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module SEDFFX1 ( SI, SE, D, CK, E, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule
module SEDFFX2 ( SI, SE, D, CK, E, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule
module SEDFFX4 ( SI, SE, D, CK, E, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule
module SEDFFXL ( SI, SE, D, CK, E, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule
module TBUFIX1 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFIX12 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFIX16 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFIX2 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFIX20 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFIX3 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFIX4 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFIX8 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFIXL ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFX1 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFX12 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFX16 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFX2 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFX20 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFX3 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFX4 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFX8 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TBUFXL ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule
module TIEHI ( Y);
    output		Y ;

endmodule
module TIELO ( Y);
    output		Y ;

endmodule
module TLATNRX1 ( D, GN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNRX2 ( D, GN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNRX4 ( D, GN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNRXL ( D, GN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNSRX1 ( D, GN, SN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNSRX2 ( D, GN, SN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNSRX4 ( D, GN, SN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNSRXL ( D, GN, SN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNSX1 ( D, GN, SN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNSX2 ( D, GN, SN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNSX4 ( D, GN, SN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNSXL ( D, GN, SN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNX1 ( D, GN, Q, QN);
    input		D ;
    input		GN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNX2 ( D, GN, Q, QN);
    input		D ;
    input		GN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNX4 ( D, GN, Q, QN);
    input		D ;
    input		GN ;
    output		Q ;
    output		QN ;

endmodule
module TLATNXL ( D, GN, Q, QN);
    input		D ;
    input		GN ;
    output		Q ;
    output		QN ;

endmodule
module TLATRX1 ( D, G, RN, Q, QN);
    input		D ;
    input		G ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATRX2 ( D, G, RN, Q, QN);
    input		D ;
    input		G ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATRX4 ( D, G, RN, Q, QN);
    input		D ;
    input		G ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATRXL ( D, G, RN, Q, QN);
    input		D ;
    input		G ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATSRX1 ( D, G, SN, RN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATSRX2 ( D, G, SN, RN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATSRX4 ( D, G, SN, RN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATSRXL ( D, G, SN, RN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule
module TLATSX1 ( D, G, SN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module TLATSX2 ( D, G, SN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module TLATSX4 ( D, G, SN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module TLATSXL ( D, G, SN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule
module TLATX1 ( D, G, Q, QN);
    input		D ;
    input		G ;
    output		Q ;
    output		QN ;

endmodule
module TLATX2 ( D, G, Q, QN);
    input		D ;
    input		G ;
    output		Q ;
    output		QN ;

endmodule
module TLATX4 ( D, G, Q, QN);
    input		D ;
    input		G ;
    output		Q ;
    output		QN ;

endmodule
module TLATXL ( D, G, Q, QN);
    input		D ;
    input		G ;
    output		Q ;
    output		QN ;

endmodule
module TTLATX1 ( D, G, OE, Q);
    input		D ;
    input		G ;
    input		OE ;
    output		Q ;

endmodule
module TTLATX2 ( D, G, OE, Q);
    input		D ;
    input		G ;
    input		OE ;
    output		Q ;

endmodule
module TTLATX4 ( D, G, OE, Q);
    input		D ;
    input		G ;
    input		OE ;
    output		Q ;

endmodule
module TTLATXL ( D, G, OE, Q);
    input		D ;
    input		G ;
    input		OE ;
    output		Q ;

endmodule
module XNOR2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module XNOR2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module XNOR2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module XNOR2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module XNOR3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module XNOR3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module XOR2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module XOR2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module XOR2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module XOR2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule
module XOR3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module XOR3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule
module PDB04DGZ ( I, OEN, PAD, C);
    input		I ;
    input		OEN ;
    inout		PAD ;
    output		C ;

endmodule
module PDIDGZ ( PAD, C);
    input		PAD ;
    output		C ;

endmodule
module PDO04CDG ( I, PAD);
    input		I ;
    output		PAD ;

endmodule
module PVDD1DGZ ( );

endmodule
module PVSS1DGZ ( );

endmodule
module PCORNERDG ( );

endmodule

# Process antenna report created by VERIFY ANTENNA.

# No Violations Found

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

NAMESCASESENSITIVE ON ;
VERSION 5.4 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO tdsp_core 
  PIN clk 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 58.1904 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 33.348 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 132.182 LAYER Metal4 ;
    ANTENNAMAXAREACAR 73.9637 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 285.101 LAYER Metal4 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 2.6544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0488 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 2.304 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 62.9328 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 240.323 LAYER Metal4 ;
    ANTENNAMAXAREACAR 64.4148 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 248.506 LAYER Metal4 ;
  END reset
  PIN as 
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 8.6744 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.1356 LAYER Metal3 ;
    ANTENNAMAXAREACAR 81.9157 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 321.926 LAYER Metal3 ;
  END as
  PIN read 
    ANTENNAPARTIALMETALAREA 3.948 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.946 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 9.3632 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.04 LAYER Metal4 ;
    ANTENNAMAXAREACAR 104.016 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 408.828 LAYER Metal4 ;
  END read
  PIN write 
    ANTENNADIFFAREA 0.924 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.6544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0488 LAYER Metal3 ;
  END write
  PIN address[7] 
    ANTENNAPARTIALMETALAREA 0.8064 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0528 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 40.4096 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 153.573 LAYER Metal4 ;
  END address[7]
  PIN address[6] 
    ANTENNAPARTIALMETALAREA 3.948 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.946 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 33.5104 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 127.454 LAYER Metal4 ;
  END address[6]
  PIN address[5] 
    ANTENNAPARTIALMETALAREA 3.7632 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2464 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 9.856 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 37.6088 LAYER Metal4 ;
  END address[5]
  PIN address[4] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 37.1392 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 140.895 LAYER Metal4 ;
  END address[4]
  PIN address[3] 
    ANTENNAPARTIALMETALAREA 0.1736 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.9927 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 20.3616 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 77.38 LAYER Metal4 ;
  END address[3]
  PIN address[2] 
    ANTENNAPARTIALMETALAREA 1.5456 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8512 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.9927 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 34.944 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 132.585 LAYER Metal4 ;
  END address[2]
  PIN address[1] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.9927 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 29.456 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 111.809 LAYER Metal4 ;
  END address[1]
  PIN address[0] 
    ANTENNAPARTIALMETALAREA 0.6216 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3532 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.6864 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 36.8032 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 139.92 LAYER Metal4 ;
  END address[0]
  PIN t_data_in[15] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.95 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.68 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9536 LAYER Metal4 ;
    ANTENNAMAXAREACAR 74.2037 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 289.095 LAYER Metal4 ;
  END t_data_in[15]
  PIN t_data_in[14] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0672 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2544 LAYER Metal3 ;
    ANTENNAMAXAREACAR 75.3444 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 290.666 LAYER Metal3 ;
  END t_data_in[14]
  PIN t_data_in[13] 
    ANTENNAPARTIALMETALAREA 0.9912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7524 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 11.2672 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.9512 LAYER Metal4 ;
    ANTENNAMAXAREACAR 68.6815 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 265.442 LAYER Metal4 ;
  END t_data_in[13]
  PIN t_data_in[12] 
    ANTENNAPARTIALMETALAREA 1.3608 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1516 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.1136 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.084 LAYER Metal4 ;
    ANTENNAMAXAREACAR 37.4148 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 147.075 LAYER Metal4 ;
  END t_data_in[12]
  PIN t_data_in[11] 
    ANTENNAPARTIALMETALAREA 5.9808 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6416 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.4272 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.2712 LAYER Metal4 ;
    ANTENNAMAXAREACAR 25.8 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 103.105 LAYER Metal4 ;
  END t_data_in[11]
  PIN t_data_in[10] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 8.736 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.6656 LAYER Metal4 ;
    ANTENNAMAXAREACAR 83.2519 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 321.975 LAYER Metal4 ;
  END t_data_in[10]
  PIN t_data_in[9] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.95 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 8.7584 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.4536 LAYER Metal4 ;
    ANTENNAMAXAREACAR 68.6296 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 265.245 LAYER Metal4 ;
  END t_data_in[9]
  PIN t_data_in[8] 
    ANTENNAPARTIALMETALAREA 1.148 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.8592 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3352 LAYER Metal4 ;
    ANTENNAMAXAREACAR 35.0296 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 138.045 LAYER Metal4 ;
  END t_data_in[8]
  PIN t_data_in[7] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.3912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3492 LAYER Metal3 ;
    ANTENNAMAXAREACAR 28.9241 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 114.931 LAYER Metal3 ;
  END t_data_in[7]
  PIN t_data_in[6] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.95 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.232 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9608 LAYER Metal4 ;
    ANTENNAMAXAREACAR 9.7 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 42.1546 LAYER Metal4 ;
  END t_data_in[6]
  PIN t_data_in[5] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.6544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0488 LAYER Metal3 ;
    ANTENNAMAXAREACAR 30.8037 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 120.673 LAYER Metal3 ;
  END t_data_in[5]
  PIN t_data_in[4] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3608 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1516 LAYER Metal3 ;
    ANTENNAMAXAREACAR 11.7481 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 48.5343 LAYER Metal3 ;
  END t_data_in[4]
  PIN t_data_in[3] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.6048 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5864 LAYER Metal4 ;
    ANTENNAMAXAREACAR 13.8481 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 57.8583 LAYER Metal4 ;
  END t_data_in[3]
  PIN t_data_in[2] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.6544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0488 LAYER Metal3 ;
    ANTENNAMAXAREACAR 16.1556 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 65.2194 LAYER Metal3 ;
  END t_data_in[2]
  PIN t_data_in[1] 
    ANTENNAPARTIALMETALAREA 1.3608 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1516 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.5456 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.148 LAYER Metal4 ;
    ANTENNAMAXAREACAR 40.3185 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 158.068 LAYER Metal4 ;
  END t_data_in[1]
  PIN t_data_in[0] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3608 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1516 LAYER Metal3 ;
    ANTENNAMAXAREACAR 10.1667 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 42.5472 LAYER Metal3 ;
  END t_data_in[0]
  PIN t_data_out[15] 
    ANTENNAPARTIALMETALAREA 0.0672 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2544 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.7845 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 11.5584 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.3504 LAYER Metal4 ;
  END t_data_out[15]
  PIN t_data_out[14] 
    ANTENNAPARTIALMETALAREA 0.6216 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3532 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.7845 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 20.9888 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 79.7544 LAYER Metal4 ;
  END t_data_out[14]
  PIN t_data_out[13] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.9184 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7736 LAYER Metal4 ;
  END t_data_out[13]
  PIN t_data_out[12] 
    ANTENNAPARTIALMETALAREA 1.148 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.9927 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 7.1456 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9416 LAYER Metal4 ;
  END t_data_out[12]
  PIN t_data_out[11] 
    ANTENNAPARTIALMETALAREA 4.1328 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6456 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 72.24 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 274.074 LAYER Metal4 ;
  END t_data_out[11]
  PIN t_data_out[10] 
    ANTENNAPARTIALMETALAREA 2.6544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0488 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 93.2288 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 353.828 LAYER Metal4 ;
  END t_data_out[10]
  PIN t_data_out[9] 
    ANTENNAPARTIALMETALAREA 0.8064 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0528 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 1.2324 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.5456 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.148 LAYER Metal4 ;
  END t_data_out[9]
  PIN t_data_out[8] 
    ANTENNAPARTIALMETALAREA 1.5456 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8512 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.7845 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 99.9712 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 379.353 LAYER Metal4 ;
  END t_data_out[8]
  PIN t_data_out[7] 
    ANTENNAPARTIALMETALAREA 1.3608 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1516 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.9927 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.3888 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5544 LAYER Metal4 ;
  END t_data_out[7]
  PIN t_data_out[6] 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 1.2324 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.7616 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.18 LAYER Metal4 ;
  END t_data_out[6]
  PIN t_data_out[5] 
    ANTENNAPARTIALMETALAREA 2.6544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0488 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 1.2324 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.0752 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3672 LAYER Metal4 ;
  END t_data_out[5]
  PIN t_data_out[4] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0672 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2544 LAYER Metal3 ;
  END t_data_out[4]
  PIN t_data_out[3] 
    ANTENNADIFFAREA 0.9927 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.9912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7524 LAYER Metal3 ;
  END t_data_out[3]
  PIN t_data_out[2] 
    ANTENNAPARTIALMETALAREA 2.4696 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3492 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 93.7216 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 355.397 LAYER Metal4 ;
  END t_data_out[2]
  PIN t_data_out[1] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 1.2324 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.7024 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7416 LAYER Metal4 ;
  END t_data_out[1]
  PIN t_data_out[0] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.9344 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7024 LAYER Metal4 ;
  END t_data_out[0]
  PIN p_read 
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 6.5632 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.44 LAYER Metal3 ;
    ANTENNAMAXAREACAR 56.9404 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 229.667 LAYER Metal3 ;
  END p_read
  PIN p_address[8] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 4.0544 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6456 LAYER Metal4 ;
  END p_address[8]
  PIN p_address[7] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.95 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 7.168 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7296 LAYER Metal4 ;
  END p_address[7]
  PIN p_address[6] 
    ANTENNAPARTIALMETALAREA 2.8392 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7484 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 11.2672 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.9512 LAYER Metal4 ;
  END p_address[6]
  PIN p_address[5] 
    ANTENNAPARTIALMETALAREA 0.8064 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0528 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 11.5808 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.1384 LAYER Metal4 ;
  END p_address[5]
  PIN p_address[4] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.024 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.448 LAYER Metal3 ;
  END p_address[4]
  PIN p_address[3] 
    ANTENNAPARTIALMETALAREA 0.9912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7524 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 16.7552 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 63.7272 LAYER Metal4 ;
  END p_address[3]
  PIN p_address[2] 
    ANTENNAPARTIALMETALAREA 0.6216 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3532 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 20.048 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 76.1928 LAYER Metal4 ;
  END p_address[2]
  PIN p_address[1] 
    ANTENNAPARTIALMETALAREA 1.3608 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1516 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 17.2032 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 65.72 LAYER Metal4 ;
  END p_address[1]
  PIN p_address[0] 
    ANTENNAPARTIALMETALAREA 3.2088 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1476 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 25.536 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 96.9688 LAYER Metal4 ;
  END p_address[0]
  PIN rom_data_in[15] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.95 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.9184 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7736 LAYER Metal4 ;
    ANTENNAMAXAREACAR 29.9222 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 118.71 LAYER Metal4 ;
  END rom_data_in[15]
  PIN rom_data_in[14] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.448 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9928 LAYER Metal4 ;
    ANTENNAMAXAREACAR 36.0407 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 141.873 LAYER Metal4 ;
  END rom_data_in[14]
  PIN rom_data_in[13] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 8.568 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.436 LAYER Metal3 ;
    ANTENNAMAXAREACAR 49.4704 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 191.34 LAYER Metal3 ;
  END rom_data_in[13]
  PIN rom_data_in[12] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
    ANTENNAMAXAREACAR 25.3333 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 99.9639 LAYER Metal3 ;
  END rom_data_in[12]
  PIN rom_data_in[11] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.2848 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6496 LAYER Metal3 ;
    ANTENNAMAXAREACAR 20.4463 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 81.463 LAYER Metal3 ;
  END rom_data_in[11]
  PIN rom_data_in[10] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER Metal3 ;
    ANTENNAMAXAREACAR 10.1667 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 42.5472 LAYER Metal3 ;
  END rom_data_in[10]
  PIN rom_data_in[9] 
    ANTENNAPARTIALMETALAREA 1.7304 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5508 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 5.4656 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.988 LAYER Metal4 ;
    ANTENNAMAXAREACAR 33.837 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 133.531 LAYER Metal4 ;
  END rom_data_in[9]
  PIN rom_data_in[8] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
    ANTENNAMAXAREACAR 13.5889 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 55.5028 LAYER Metal3 ;
  END rom_data_in[8]
  PIN rom_data_in[7] 
    ANTENNAPARTIALMETALAREA 9.6768 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.6336 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.1136 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.084 LAYER Metal4 ;
    ANTENNAMAXAREACAR 18.4111 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 75.1324 LAYER Metal4 ;
  END rom_data_in[7]
  PIN rom_data_in[6] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.448 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9928 LAYER Metal4 ;
    ANTENNAMAXAREACAR 69.9259 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 270.153 LAYER Metal4 ;
  END rom_data_in[6]
  PIN rom_data_in[5] 
    ANTENNAPARTIALMETALAREA 1.7304 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5508 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.6432 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3032 LAYER Metal4 ;
    ANTENNAMAXAREACAR 19.4611 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 79.1074 LAYER Metal4 ;
  END rom_data_in[5]
  PIN rom_data_in[4] 
    ANTENNAPARTIALMETALAREA 3.7632 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2464 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.9184 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7736 LAYER Metal4 ;
    ANTENNAMAXAREACAR 59.6074 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 231.09 LAYER Metal4 ;
  END rom_data_in[4]
  PIN rom_data_in[3] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.896 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9856 LAYER Metal4 ;
    ANTENNAMAXAREACAR 58.9333 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 231.286 LAYER Metal4 ;
  END rom_data_in[3]
  PIN rom_data_in[2] 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 15.5008 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 58.9784 LAYER Metal4 ;
    ANTENNAMAXAREACAR 125.381 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 480.092 LAYER Metal4 ;
  END rom_data_in[2]
  PIN rom_data_in[1] 
    ANTENNAPARTIALMETALAREA 3.7632 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2464 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.8592 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3352 LAYER Metal4 ;
    ANTENNAMAXAREACAR 47.6296 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 185.745 LAYER Metal4 ;
  END rom_data_in[1]
  PIN rom_data_in[0] 
    ANTENNAPARTIALMETALAREA 0.0672 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2544 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 12.9696 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 49.6928 LAYER Metal4 ;
    ANTENNAMAXAREACAR 125.511 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 483.331 LAYER Metal4 ;
  END rom_data_in[0]
  PIN bus_grant 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 1.4331 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 37.8112 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 144.923 LAYER Metal4 ;
    ANTENNAMAXAREACAR 48.5452 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 187.315 LAYER Metal4 ;
  END bus_grant
  PIN bus_request 
    ANTENNAPARTIALMETALAREA 1.176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.6846 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 39.4016 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 150.647 LAYER Metal4 ;
    ANTENNAMAXAREACAR 130.185 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 499.607 LAYER Metal4 ;
  END bus_request
  PIN port_as 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.1008 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 14.6944 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 56.2224 LAYER Metal4 ;
    ANTENNAMAXAREACAR 458.778 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 1754.68 LAYER Metal4 ;
  END port_as
  PIN port_address[2] 
    ANTENNAPARTIALMETALAREA 4.1328 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6456 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 10.1472 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.008 LAYER Metal4 ;
  END port_address[2]
  PIN port_address[1] 
    ANTENNAPARTIALMETALAREA 4.1328 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6456 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.6864 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.6048 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5864 LAYER Metal4 ;
  END port_address[1]
  PIN port_address[0] 
    ANTENNAPARTIALMETALAREA 3.948 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.946 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.6864 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.0752 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3672 LAYER Metal4 ;
  END port_address[0]
  PIN port_pad_data_in[15] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.6216 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3532 LAYER Metal3 ;
    ANTENNAMAXAREACAR 11.9556 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 49.3194 LAYER Metal3 ;
  END port_pad_data_in[15]
  PIN port_pad_data_in[14] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 16.5144 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.5188 LAYER Metal3 ;
    ANTENNAMAXAREACAR 86.9852 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 333.36 LAYER Metal3 ;
  END port_pad_data_in[14]
  PIN port_pad_data_in[13] 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 18.7488 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 71.868 LAYER Metal4 ;
    ANTENNAMAXAREACAR 146.9 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 565.677 LAYER Metal4 ;
  END port_pad_data_in[13]
  PIN port_pad_data_in[12] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.7616 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.18 LAYER Metal4 ;
    ANTENNAMAXAREACAR 77.2111 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 299.106 LAYER Metal4 ;
  END port_pad_data_in[12]
  PIN port_pad_data_in[11] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.652 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5508 LAYER Metal3 ;
    ANTENNAMAXAREACAR 23.9852 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 96.2343 LAYER Metal3 ;
  END port_pad_data_in[11]
  PIN port_pad_data_in[10] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.4696 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3492 LAYER Metal3 ;
    ANTENNAMAXAREACAR 69.563 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 271.527 LAYER Metal3 ;
  END port_pad_data_in[10]
  PIN port_pad_data_in[9] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAMAXAREACAR 38.4519 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 151.001 LAYER Metal3 ;
  END port_pad_data_in[9]
  PIN port_pad_data_in[8] 
    ANTENNAPARTIALMETALAREA 0.9912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7524 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.7408 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4584 LAYER Metal4 ;
    ANTENNAMAXAREACAR 50.1444 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 196.64 LAYER Metal4 ;
  END port_pad_data_in[8]
  PIN port_pad_data_in[7] 
    ANTENNAPARTIALMETALAREA 2.3912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3492 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.7616 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.18 LAYER Metal4 ;
    ANTENNAMAXAREACAR 13.6407 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 59.8213 LAYER Metal4 ;
  END port_pad_data_in[7]
  PIN port_pad_data_in[6] 
    ANTENNAPARTIALMETALAREA 2.6544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0488 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.1136 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.084 LAYER Metal4 ;
    ANTENNAMAXAREACAR 30.8815 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 122.342 LAYER Metal4 ;
  END port_pad_data_in[6]
  PIN port_pad_data_in[5] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER Metal3 ;
    ANTENNAMAXAREACAR 42.1074 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 163.466 LAYER Metal3 ;
  END port_pad_data_in[5]
  PIN port_pad_data_in[4] 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.232 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9608 LAYER Metal4 ;
    ANTENNAMAXAREACAR 53.0481 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 206.258 LAYER Metal4 ;
  END port_pad_data_in[4]
  PIN port_pad_data_in[3] 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.2088 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1476 LAYER Metal3 ;
    ANTENNAMAXAREACAR 58.0519 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 223.827 LAYER Metal3 ;
  END port_pad_data_in[3]
  PIN port_pad_data_in[2] 
    ANTENNAPARTIALMETALAREA 0.9912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7524 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 9.0496 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.8528 LAYER Metal4 ;
    ANTENNAMAXAREACAR 59.0889 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 230.501 LAYER Metal4 ;
  END port_pad_data_in[2]
  PIN port_pad_data_in[1] 
    ANTENNAPARTIALMETALAREA 12.4488 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.1276 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.8304 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.688 LAYER Metal4 ;
    ANTENNAMAXAREACAR 42.0296 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 168.668 LAYER Metal4 ;
  END port_pad_data_in[1]
  PIN port_pad_data_in[0] 
    ANTENNAPARTIALMETALAREA 3.3936 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.8472 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.216 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.1136 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.084 LAYER Metal4 ;
    ANTENNAMAXAREACAR 37.4148 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 147.075 LAYER Metal4 ;
  END port_pad_data_in[0]
  PIN port_pad_data_out[15] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0672 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2544 LAYER Metal3 ;
  END port_pad_data_out[15]
  PIN port_pad_data_out[14] 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 24.752 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 94.0008 LAYER Metal4 ;
  END port_pad_data_out[14]
  PIN port_pad_data_out[13] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 31.9592 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 121.285 LAYER Metal3 ;
  END port_pad_data_out[13]
  PIN port_pad_data_out[12] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER Metal3 ;
  END port_pad_data_out[12]
  PIN port_pad_data_out[11] 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.8 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8968 LAYER Metal4 ;
  END port_pad_data_out[11]
  PIN port_pad_data_out[10] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.8976 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.052 LAYER Metal4 ;
  END port_pad_data_out[10]
  PIN port_pad_data_out[9] 
    ANTENNAPARTIALMETALAREA 0.9912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7524 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.6432 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3032 LAYER Metal4 ;
  END port_pad_data_out[9]
  PIN port_pad_data_out[8] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0672 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2544 LAYER Metal3 ;
  END port_pad_data_out[8]
  PIN port_pad_data_out[7] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0672 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2544 LAYER Metal3 ;
  END port_pad_data_out[7]
  PIN port_pad_data_out[6] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
  END port_pad_data_out[6]
  PIN port_pad_data_out[5] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
  END port_pad_data_out[5]
  PIN port_pad_data_out[4] 
    ANTENNADIFFAREA 0.5544 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.9912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7524 LAYER Metal3 ;
  END port_pad_data_out[4]
  PIN port_pad_data_out[3] 
    ANTENNAPARTIALMETALAREA 4.1328 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6456 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.0752 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3672 LAYER Metal4 ;
  END port_pad_data_out[3]
  PIN port_pad_data_out[2] 
    ANTENNAPARTIALMETALAREA 3.948 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.946 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 6.384 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.7616 LAYER Metal4 ;
  END port_pad_data_out[2]
  PIN port_pad_data_out[1] 
    ANTENNAPARTIALMETALAREA 5.0568 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1436 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.7408 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4584 LAYER Metal4 ;
  END port_pad_data_out[1]
  PIN port_pad_data_out[0] 
    ANTENNAPARTIALMETALAREA 1.176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNADIFFAREA 0.6864 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.2704 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6776 LAYER Metal4 ;
  END port_pad_data_out[0]
  PIN bio 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.108 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.2912 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3992 LAYER Metal4 ;
    ANTENNAMAXAREACAR 60.2593 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 245.272 LAYER Metal4 ;
  END bio
  PIN int 
    ANTENNAGATEAREA 0.108 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 1.176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER Metal3 ;
    ANTENNAMAXAREACAR 30.4963 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 127.102 LAYER Metal3 ;
  END int
  PIN scan_en 
    ANTENNAPARTIALMETALAREA 4.3176 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 68.3928 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 69.8432 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 277.466 LAYER Metal4 ;
    ANTENNAMAXAREACAR 78.4354 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 304.301 LAYER Metal4 ;
  END scan_en
  PIN BG_scan_in 
  END BG_scan_in
  PIN BG_scan_out 
    ANTENNAPARTIALMETALAREA 62.2664 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 236.02 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.5544 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.8368 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5472 LAYER Metal4 ;
    ANTENNAMAXAREACAR 51.8619 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 211.387 LAYER Metal4 ;
  END BG_scan_out
  PIN SPCASCAN_N1_p_data_out_13_ 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 7.8288 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.6376 LAYER Metal3 ;
    ANTENNAMAXAREACAR 39.6965 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 154.044 LAYER Metal3 ;
#    ANTENNAGATEAREA 0.216 LAYER Via34 ; 
#    ANTENNADIFFAREA 0.924 LAYER Via34 ; 
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAMAXCUTCAR 0.938889 LAYER Via34 ;
    ANTENNAGATEAREA 0.792 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 87.6064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 332.246 LAYER Metal4 ;
    ANTENNAMAXAREACAR 165.816 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 631.025 LAYER Metal4 ;
  END SPCASCAN_N1_p_data_out_13_
  PIN SPCASCAN_N2_low_mag_8_ 
    ANTENNAPARTIALMETALAREA 1.9152 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2504 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.2912 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3992 LAYER Metal4 ;
    ANTENNAMAXAREACAR 75.9095 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 299.188 LAYER Metal4 ;
  END SPCASCAN_N2_low_mag_8_
  PIN SPCASCAN_N3_port_data_out_0_ 
    ANTENNAGATEAREA 0.6153 LAYER Metal3 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 69.9776 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 266.102 LAYER Metal3 ;
    ANTENNAMAXAREACAR 144.095 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 551.997 LAYER Metal3 ;
  END SPCASCAN_N3_port_data_out_0_
  PIN SPCASCAN_N4_low_mag_3_ 
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.024 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.448 LAYER Metal3 ;
    ANTENNAMAXAREACAR 39.5268 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 159.164 LAYER Metal3 ;
  END SPCASCAN_N4_low_mag_3_
  PIN SPCASCAN_N5_port_data_out_1_ 
    ANTENNAPARTIALMETALAREA 0.9912 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7524 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.6153 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 134.316 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 509.669 LAYER Metal4 ;
    ANTENNAMAXAREACAR 246.427 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 938.596 LAYER Metal4 ;
  END SPCASCAN_N5_port_data_out_1_
  PIN FE_PT1_ 
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.2848 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6496 LAYER Metal3 ;
    ANTENNAMAXAREACAR 81.1595 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 319.063 LAYER Metal3 ;
  END FE_PT1_
  PIN SPCASCAN_N22_data_out_0_ 
    ANTENNAPARTIALMETALAREA 0.0672 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2544 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.4068 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.4416 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1336 LAYER Metal4 ;
    ANTENNAMAXAREACAR 35.1985 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 139.204 LAYER Metal4 ;
  END SPCASCAN_N22_data_out_0_
  PIN SPCASCAN_N24_t_sel_7 
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.7632 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2464 LAYER Metal3 ;
    ANTENNAMAXAREACAR 47.6503 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 189.917 LAYER Metal3 ;
  END SPCASCAN_N24_t_sel_7
  PIN SPCASCAN_N25_data_out_12_ 
    ANTENNAGATEAREA 0.216 LAYER Metal3 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 4.2392 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3452 LAYER Metal3 ;
    ANTENNAMAXAREACAR 31.3873 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 123.961 LAYER Metal3 ;
#    ANTENNAGATEAREA 0.216 LAYER Via34 ; 
#    ANTENNADIFFAREA 0.924 LAYER Via34 ; 
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAMAXCUTCAR 1.25185 LAYER Via34 ;
    ANTENNAGATEAREA 0.4068 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 7.0336 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 26.924 LAYER Metal4 ;
    ANTENNAMAXAREACAR 48.6773 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 190.146 LAYER Metal4 ;
  END SPCASCAN_N25_data_out_12_
  PIN SPCASCAN_N26_spi_sr_0_ 
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.5784 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.5468 LAYER Metal3 ;
    ANTENNAMAXAREACAR 35.1397 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 143.501 LAYER Metal3 ;
  END SPCASCAN_N26_spi_sr_0_
  PIN SPCASCAN_N27_port_data_out_11_ 
    ANTENNAPARTIALMETALAREA 0.8064 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0528 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.6153 LAYER Metal4 ; 
    ANTENNADIFFAREA 0.924 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 4.2672 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.3416 LAYER Metal4 ;
    ANTENNAMAXAREACAR 26.9502 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 106.523 LAYER Metal4 ;
  END SPCASCAN_N27_port_data_out_11_
  PIN n_7862 
    ANTENNAPARTIALMETALAREA 24.752 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 94.0008 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAGATEAREA 0.1008 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.0752 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3672 LAYER Metal4 ;
    ANTENNAMAXAREACAR 17.2778 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 77.3968 LAYER Metal4 ;
  END n_7862
##  PIN VDD 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD
#  PIN VDD.extra1 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra1
#  PIN VDD.extra2 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra2
#  PIN VDD.extra3 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra3
#  PIN VDD.extra4 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra4
#  PIN VDD.extra5 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra5
#  PIN VDD.extra6 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra6
#  PIN VDD.extra7 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra7
#  PIN VDD.extra8 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra8
#  PIN VDD.extra9 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra9
#  PIN VDD.extra10 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra10
#  PIN VDD.extra11 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra11
#  PIN VDD.extra12 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra12
#  PIN VDD.extra13 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra13
#  PIN VDD.extra14 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra14
#  PIN VDD.extra15 
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra15
#  PIN VDD.extra16 
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra16
#  PIN VDD.extra17 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra17
#  PIN VDD.extra18 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra18
#  PIN VDD.extra19 
#    ANTENNAPARTIALMETALAREA 280.432 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 371.572 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra19
#  PIN VDD.extra20 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra20
#  PIN VDD.extra21 
#    ANTENNAPARTIALMETALAREA 280.432 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 371.572 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra21
#  PIN VDD.extra22 
#    ANTENNAPARTIALMETALAREA 280.432 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 371.572 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra22
#  PIN VDD.extra23 
#    ANTENNAPARTIALMETALAREA 253.024 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 335.257 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra23
#  PIN VDD.extra24 
#    ANTENNAPARTIALMETALAREA 280.432 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 371.572 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra24
#  PIN VDD.extra25 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra25
#  PIN VDD.extra26 
#    ANTENNAPARTIALMETALAREA 258.304 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 342.253 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra26
#  PIN VDD.extra27 
#    ANTENNAPARTIALMETALAREA 258.304 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 342.253 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra27
#  PIN VDD.extra28 
#    ANTENNAPARTIALMETALAREA 258.304 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 342.253 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra28
#  PIN VDD.extra29 
#    ANTENNAPARTIALMETALAREA 253.024 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 335.257 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra29
#  PIN VDD.extra30 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra30
#  PIN VDD.extra31 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra31
#  PIN VDD.extra32 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra32
#  PIN VDD.extra33 
#    ANTENNAPARTIALMETALAREA 280.432 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 371.572 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra33
#  PIN VDD.extra34 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra34
#  PIN VDD.extra35 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra35
#  PIN VDD.extra36 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra36
#  PIN VDD.extra37 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra37
#  PIN VDD.extra38 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra38
#  PIN VDD.extra39 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra39
#  PIN VDD.extra40 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra40
#  PIN VDD.extra41 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra41
#  PIN VDD.extra42 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra42
#  PIN VDD.extra43 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra43
#  PIN VDD.extra44 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra44
#  PIN VDD.extra45 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra45
#  PIN VDD.extra46 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra46
#  PIN VDD.extra47 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra47
#  PIN VDD.extra48 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra48
#  PIN VDD.extra49 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra49
#  PIN VDD.extra50 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra50
#  PIN VDD.extra51 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra51
#  PIN VDD.extra52 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra52
#  PIN VDD.extra53 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra53
#  PIN VDD.extra54 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra54
#  PIN VDD.extra55 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra55
#  PIN VDD.extra56 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra56
#  PIN VDD.extra57 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra57
#  PIN VDD.extra58 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra58
#  PIN VDD.extra59 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra59
#  PIN VDD.extra60 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra60
#  PIN VDD.extra61 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra61
#  PIN VDD.extra62 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6382 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1403.44 LAYER Metal4 ;
#  END VDD.extra62
#  PIN VSS 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS
#  PIN VSS.extra1 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra1
#  PIN VSS.extra2 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra2
#  PIN VSS.extra3 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra3
#  PIN VSS.extra4 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra4
#  PIN VSS.extra5 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra5
#  PIN VSS.extra6 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra6
#  PIN VSS.extra7 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra7
#  PIN VSS.extra8 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra8
#  PIN VSS.extra9 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra9
#  PIN VSS.extra10 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra10
#  PIN VSS.extra11 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra11
#  PIN VSS.extra12 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra12
#  PIN VSS.extra13 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra13
#  PIN VSS.extra14 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra14
#  PIN VSS.extra15 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra15
#  PIN VSS.extra16 
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra16
#  PIN VSS.extra17 
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra17
#  PIN VSS.extra18 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra18
#  PIN VSS.extra19 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra19
#  PIN VSS.extra20 
#    ANTENNAPARTIALMETALAREA 287.312 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 380.688 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra20
#  PIN VSS.extra21 
#    ANTENNAPARTIALMETALAREA 287.312 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 380.688 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra21
#  PIN VSS.extra22 
#    ANTENNAPARTIALMETALAREA 287.312 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 380.688 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra22
#  PIN VSS.extra23 
#    ANTENNAPARTIALMETALAREA 258.304 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 342.253 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra23
#  PIN VSS.extra24 
#    ANTENNAPARTIALMETALAREA 287.312 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 380.688 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra24
#  PIN VSS.extra25 
#    ANTENNAPARTIALMETALAREA 253.024 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 335.257 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra25
#  PIN VSS.extra26 
#    ANTENNAPARTIALMETALAREA 287.312 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 380.688 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra26
#  PIN VSS.extra27 
#    ANTENNAPARTIALMETALAREA 258.304 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 342.253 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra27
#  PIN VSS.extra28 
#    ANTENNAPARTIALMETALAREA 258.304 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 342.253 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra28
#  PIN VSS.extra29 
#    ANTENNAPARTIALMETALAREA 253.552 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 335.956 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra29
#  PIN VSS.extra30 
#    ANTENNAPARTIALMETALAREA 287.312 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 380.688 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 14.4 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 21.624 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra30
#  PIN VSS.extra31 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra31
#  PIN VSS.extra32 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra32
#  PIN VSS.extra33 
#    ANTENNAPARTIALMETALAREA 255.664 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 338.755 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra33
#  PIN VSS.extra34 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra34
#  PIN VSS.extra35 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra35
#  PIN VSS.extra36 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra36
#  PIN VSS.extra37 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra37
#  PIN VSS.extra38 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra38
#  PIN VSS.extra39 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra39
#  PIN VSS.extra40 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra40
#  PIN VSS.extra41 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra41
#  PIN VSS.extra42 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra42
#  PIN VSS.extra43 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra43
#  PIN VSS.extra44 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra44
#  PIN VSS.extra45 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra45
#  PIN VSS.extra46 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra46
#  PIN VSS.extra47 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra47
#  PIN VSS.extra48 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra48
#  PIN VSS.extra49 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra49
#  PIN VSS.extra50 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra50
#  PIN VSS.extra51 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra51
#  PIN VSS.extra52 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra52
#  PIN VSS.extra53 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra53
#  PIN VSS.extra54 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra54
#  PIN VSS.extra55 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra55
#  PIN VSS.extra56 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra56
#  PIN VSS.extra57 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra57
#  PIN VSS.extra58 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra58
#  PIN VSS.extra59 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra59
#  PIN VSS.extra60 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra60
#  PIN VSS.extra61 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra61
#  PIN VSS.extra62 
#    ANTENNAPARTIALMETALAREA 354.4 LAYER Metal1 ;
#    ANTENNAPARTIALMETALSIDEAREA 469.58 LAYER Metal1 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal2 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal2 ;
#    ANTENNAPARTIALMETALAREA 8 LAYER Metal3 ;
#    ANTENNAPARTIALMETALSIDEAREA 12.296 LAYER Metal3 ;
#    ANTENNAPARTIALMETALAREA 6388.4 LAYER Metal4 ;
#    ANTENNAPARTIALMETALSIDEAREA 1412.77 LAYER Metal4 ;
#  END VSS.extra62
END tdsp_core

END LIBRARY

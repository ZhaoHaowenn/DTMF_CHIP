
module ADDFHX1 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule

module ADDFHX2 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule

module ADDFHX4 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule

module ADDFHXL ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule

module ADDFX1 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule

module ADDFX2 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule

module ADDFX4 ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule

module ADDFXL ( A, B, CI, S, CO);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CO ;

endmodule

module ADDHX1 ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule

module ADDHX2 ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule

module ADDHX4 ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule

module ADDHXL ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule

module AFCSHCINX2 ( CS, A, B, CI0N, CI1N, S, CO0, CO1);
    input		CS ;
    input		A ;
    input		B ;
    input		CI0N ;
    input		CI1N ;
    output		S ;
    output		CO0 ;
    output		CO1 ;

endmodule

module AFCSHCINX4 ( CS, A, B, CI0N, CI1N, S, CO0, CO1);
    input		CS ;
    input		A ;
    input		B ;
    input		CI0N ;
    input		CI1N ;
    output		S ;
    output		CO0 ;
    output		CO1 ;

endmodule

module AFCSHCONX2 ( CS, A, B, CI0, CI1, S, CO0N, CO1N);
    input		CS ;
    input		A ;
    input		B ;
    input		CI0 ;
    input		CI1 ;
    output		S ;
    output		CO0N ;
    output		CO1N ;

endmodule

module AFCSHCONX4 ( CS, A, B, CI0, CI1, S, CO0N, CO1N);
    input		CS ;
    input		A ;
    input		B ;
    input		CI0 ;
    input		CI1 ;
    output		S ;
    output		CO0N ;
    output		CO1N ;

endmodule

module AFHCINX2 ( A, B, CIN, S, CO);
    input		A ;
    input		B ;
    input		CIN ;
    output		S ;
    output		CO ;

endmodule

module AFHCINX4 ( A, B, CIN, S, CO);
    input		A ;
    input		B ;
    input		CIN ;
    output		S ;
    output		CO ;

endmodule

module AFHCONX2 ( A, B, CI, S, CON);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CON ;

endmodule

module AFHCONX4 ( A, B, CI, S, CON);
    input		A ;
    input		B ;
    input		CI ;
    output		S ;
    output		CON ;

endmodule

module AHHCINX2 ( A, CIN, S, CO);
    input		A ;
    input		CIN ;
    output		S ;
    output		CO ;

endmodule

module AHHCINX4 ( A, CIN, S, CO);
    input		A ;
    input		CIN ;
    output		S ;
    output		CO ;

endmodule

module AHHCONX2 ( A, CI, S, CON);
    input		A ;
    input		CI ;
    output		S ;
    output		CON ;

endmodule

module AHHCONX4 ( A, CI, S, CON);
    input		A ;
    input		CI ;
    output		S ;
    output		CON ;

endmodule

module AND2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module AND2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module AND2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module AND2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module AND3X1 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module AND3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module AND3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module AND3XL ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module AND4X1 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module AND4X2 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module AND4X4 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module AND4XL ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module AOI211X1 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule

module AOI211X2 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule

module AOI211X4 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule

module AOI211XL ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule

module AOI21X1 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule

module AOI21X2 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule

module AOI21X4 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule

module AOI21XL ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule

module AOI221X1 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule

module AOI221X2 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule

module AOI221X4 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule

module AOI221XL ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule

module AOI222X1 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule

module AOI222X2 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule

module AOI222X4 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule

module AOI222XL ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule

module AOI22X1 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI22X2 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI22X4 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI22XL ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI2BB1X1 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule

module AOI2BB1X2 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule

module AOI2BB1X4 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule

module AOI2BB1XL ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule

module AOI2BB2X1 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI2BB2X2 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI2BB2X4 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI2BB2XL ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI31X1 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule

module AOI31X2 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule

module AOI31X4 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule

module AOI31XL ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule

module AOI32X1 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI32X2 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI32X4 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI32XL ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module AOI33X1 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule

module AOI33X2 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule

module AOI33X4 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule

module AOI33XL ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule

module BENCX1 ( M2, M1, M0, A, S, X2);
    input		M2 ;
    input		M1 ;
    input		M0 ;
    output		A ;
    output		S ;
    output		X2 ;

endmodule

module BENCX2 ( M2, M1, M0, A, S, X2);
    input		M2 ;
    input		M1 ;
    input		M0 ;
    output		A ;
    output		S ;
    output		X2 ;

endmodule

module BENCX4 ( M2, M1, M0, A, S, X2);
    input		M2 ;
    input		M1 ;
    input		M0 ;
    output		A ;
    output		S ;
    output		X2 ;

endmodule

module BMXX1 ( X2, M0, A, S, M1, PP);
    input		X2 ;
    input		M0 ;
    input		A ;
    input		S ;
    input		M1 ;
    output		PP ;

endmodule

module BUFX1 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module BUFX12 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module BUFX16 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module BUFX2 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module BUFX20 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module BUFX3 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module BUFX4 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module BUFX8 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module BUFXL ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFX1 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFX12 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFX16 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFX2 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFX20 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFX3 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFX4 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFX8 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKBUFXL ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVX1 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVX12 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVX16 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVX2 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVX20 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVX3 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVX4 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVX8 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CLKINVXL ( A, Y);
    input		A ;
    output		Y ;

endmodule

module CMPR22X1 ( A, B, S, CO);
    input		A ;
    input		B ;
    output		S ;
    output		CO ;

endmodule

module CMPR32X1 ( A, B, C, S, CO);
    input		A ;
    input		B ;
    input		C ;
    output		S ;
    output		CO ;

endmodule

module CMPR42X1 ( A, B, C, D, ICI, S, ICO, CO);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    input		ICI ;
    output		S ;
    output		ICO ;
    output		CO ;

endmodule

module CMPR42X2 ( A, B, C, D, ICI, S, ICO, CO);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    input		ICI ;
    output		S ;
    output		ICO ;
    output		CO ;

endmodule

module DFFHQX1 ( D, CK, Q);
    input		D ;
    input		CK ;
    output		Q ;

endmodule

module DFFHQX2 ( D, CK, Q);
    input		D ;
    input		CK ;
    output		Q ;

endmodule

module DFFHQX4 ( D, CK, Q);
    input		D ;
    input		CK ;
    output		Q ;

endmodule

module DFFHQXL ( D, CK, Q);
    input		D ;
    input		CK ;
    output		Q ;

endmodule

module DFFNRX1 ( D, CKN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNRX2 ( D, CKN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNRX4 ( D, CKN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNRXL ( D, CKN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNSRX1 ( D, CKN, SN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNSRX2 ( D, CKN, SN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNSRX4 ( D, CKN, SN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNSRXL ( D, CKN, SN, RN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNSX1 ( D, CKN, SN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNSX2 ( D, CKN, SN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNSX4 ( D, CKN, SN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNSXL ( D, CKN, SN, Q, QN);
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNX1 ( D, CKN, Q, QN);
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNX2 ( D, CKN, Q, QN);
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNX4 ( D, CKN, Q, QN);
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule

module DFFNXL ( D, CKN, Q, QN);
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule

module DFFRHQX1 ( D, CK, RN, Q);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule

module DFFRHQX2 ( D, CK, RN, Q);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule

module DFFRHQX4 ( D, CK, RN, Q);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule

module DFFRHQXL ( D, CK, RN, Q);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule

module DFFRX1 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFRX2 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFRX4 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFRXL ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFSHQX1 ( D, CK, SN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule

module DFFSHQX2 ( D, CK, SN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule

module DFFSHQX4 ( D, CK, SN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule

module DFFSHQXL ( D, CK, SN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule

module DFFSRHQX1 ( D, CK, SN, RN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule

module DFFSRHQX2 ( D, CK, SN, RN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule

module DFFSRHQX4 ( D, CK, SN, RN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule

module DFFSRHQXL ( D, CK, SN, RN, Q);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule

module DFFSRX1 ( D, CK, SN, RN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFSRX2 ( D, CK, SN, RN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFSRX4 ( D, CK, SN, RN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFSRXL ( D, CK, SN, RN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFSX1 ( D, CK, SN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module DFFSX2 ( D, CK, SN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module DFFSX4 ( D, CK, SN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module DFFSXL ( D, CK, SN, Q, QN);
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module DFFTRX1 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFTRX2 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFTRX4 ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFTRXL ( D, CK, RN, Q, QN);
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module DFFX1 ( D, CK, Q, QN);
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module DFFX2 ( D, CK, Q, QN);
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module DFFX4 ( D, CK, Q, QN);
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module DFFXL ( D, CK, Q, QN);
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module DLY1X1 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module DLY2X1 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module DLY3X1 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module DLY4X1 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module EDFFTRX1 ( D, CK, E, RN, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module EDFFTRX2 ( D, CK, E, RN, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module EDFFTRX4 ( D, CK, E, RN, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module EDFFTRXL ( D, CK, E, RN, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module EDFFX1 ( D, CK, E, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule

module EDFFX2 ( D, CK, E, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule

module EDFFX4 ( D, CK, E, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule

module EDFFXL ( D, CK, E, Q, QN);
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule

module HOLDX1 ( Y);
    inout		Y ;

endmodule

module INVX1 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module INVX12 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module INVX16 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module INVX2 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module INVX20 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module INVX3 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module INVX4 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module INVX8 ( A, Y);
    input		A ;
    output		Y ;

endmodule

module INVXL ( A, Y);
    input		A ;
    output		Y ;

endmodule

module JKFFRX1 ( J, K, CK, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFRX2 ( J, K, CK, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFRX4 ( J, K, CK, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFRXL ( J, K, CK, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFSRX1 ( J, K, CK, SN, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFSRX2 ( J, K, CK, SN, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFSRX4 ( J, K, CK, SN, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFSRXL ( J, K, CK, SN, RN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFSX1 ( J, K, CK, SN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFSX2 ( J, K, CK, SN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFSX4 ( J, K, CK, SN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFSXL ( J, K, CK, SN, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module JKFFX1 ( J, K, CK, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module JKFFX2 ( J, K, CK, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module JKFFX4 ( J, K, CK, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module JKFFXL ( J, K, CK, Q, QN);
    input		J ;
    input		K ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module MX2X1 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MX2X2 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MX2X4 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MX2XL ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MX4X1 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MX4X2 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MX4X4 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MX4XL ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MXI2X1 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MXI2X2 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MXI2X4 ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MXI2XL ( S0, B, A, Y);
    input		S0 ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MXI4X1 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MXI4X2 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MXI4X4 ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module MXI4XL ( S1, S0, D, C, B, A, Y);
    input		S1 ;
    input		S0 ;
    input		D ;
    input		C ;
    input		B ;
    input		A ;
    output		Y ;

endmodule

module NAND2BX1 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule

module NAND2BX2 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule

module NAND2BX4 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule

module NAND2BXL ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule

module NAND2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module NAND2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module NAND2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module NAND2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module NAND3BX1 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NAND3BX2 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NAND3BX4 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NAND3BXL ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NAND3X1 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NAND3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NAND3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NAND3XL ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NAND4BBX1 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4BBX2 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4BBX4 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4BBXL ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4BX1 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4BX2 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4BX4 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4BXL ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4X1 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4X2 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4X4 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NAND4XL ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR2BX1 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule

module NOR2BX2 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule

module NOR2BX4 ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule

module NOR2BXL ( AN, B, Y);
    input		AN ;
    input		B ;
    output		Y ;

endmodule

module NOR2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module NOR2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module NOR2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module NOR2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module NOR3BX1 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NOR3BX2 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NOR3BX4 ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NOR3BXL ( AN, B, C, Y);
    input		AN ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NOR3X1 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NOR3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NOR3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NOR3XL ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module NOR4BBX1 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4BBX2 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4BBX4 ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4BBXL ( AN, BN, C, D, Y);
    input		AN ;
    input		BN ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4BX1 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4BX2 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4BX4 ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4BXL ( AN, B, C, D, Y);
    input		AN ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4X1 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4X2 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4X4 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module NOR4XL ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module OAI211X1 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule

module OAI211X2 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule

module OAI211X4 ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule

module OAI211XL ( A0, A1, B0, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		C0 ;
    output		Y ;

endmodule

module OAI21X1 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule

module OAI21X2 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule

module OAI21X4 ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule

module OAI21XL ( A0, A1, B0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    output		Y ;

endmodule

module OAI221X1 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule

module OAI221X2 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule

module OAI221X4 ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule

module OAI221XL ( A0, A1, B0, B1, C0, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    output		Y ;

endmodule

module OAI222X1 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule

module OAI222X2 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule

module OAI222X4 ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule

module OAI222XL ( A0, A1, B0, B1, C0, C1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    input		C0 ;
    input		C1 ;
    output		Y ;

endmodule

module OAI22X1 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI22X2 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI22X4 ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI22XL ( A0, A1, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI2BB1X1 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule

module OAI2BB1X2 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule

module OAI2BB1X4 ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule

module OAI2BB1XL ( A0N, A1N, B0, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    output		Y ;

endmodule

module OAI2BB2X1 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI2BB2X2 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI2BB2X4 ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI2BB2XL ( A0N, A1N, B0, B1, Y);
    input		A0N ;
    input		A1N ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI31X1 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule

module OAI31X2 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule

module OAI31X4 ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule

module OAI31XL ( A0, A1, A2, B0, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    output		Y ;

endmodule

module OAI32X1 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI32X2 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI32X4 ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI32XL ( A0, A1, A2, B0, B1, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    output		Y ;

endmodule

module OAI33X1 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule

module OAI33X2 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule

module OAI33X4 ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule

module OAI33XL ( A0, A1, A2, B0, B1, B2, Y);
    input		A0 ;
    input		A1 ;
    input		A2 ;
    input		B0 ;
    input		B1 ;
    input		B2 ;
    output		Y ;

endmodule

module OR2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module OR2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module OR2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module OR2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module OR3X1 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module OR3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module OR3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module OR3XL ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module OR4X1 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module OR4X2 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module OR4X4 ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module OR4XL ( A, B, C, D, Y);
    input		A ;
    input		B ;
    input		C ;
    input		D ;
    output		Y ;

endmodule

module RF1R1WX2 ( WW, WB, RW, RWN, RB);
    input		WW ;
    input		WB ;
    input		RW ;
    input		RWN ;
    output		RB ;

endmodule

module RF2R1WX2 ( WB, WW, R1W, R2W, R1B, R2B);
    input		WB ;
    input		WW ;
    input		R1W ;
    input		R2W ;
    output		R1B ;
    output		R2B ;

endmodule

module RFRDX1 ( RB, BRB);
    input		RB ;
    output		BRB ;

endmodule

module RFRDX2 ( RB, BRB);
    input		RB ;
    output		BRB ;

endmodule

module RFRDX4 ( RB, BRB);
    input		RB ;
    output		BRB ;

endmodule

module SDFFHQX1 ( SI, SE, D, CK, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;

endmodule

module SDFFHQX2 ( SI, SE, D, CK, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;

endmodule

module SDFFHQX4 ( SI, SE, D, CK, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;

endmodule

module SDFFHQXL ( SI, SE, D, CK, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;

endmodule

module SDFFNRX1 ( SI, SE, D, CKN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNRX2 ( SI, SE, D, CKN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNRX4 ( SI, SE, D, CKN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNRXL ( SI, SE, D, CKN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNSRX1 ( SI, SE, D, CKN, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNSRX2 ( SI, SE, D, CKN, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNSRX4 ( SI, SE, D, CKN, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNSRXL ( SI, SE, D, CKN, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNSX1 ( SI, SE, D, CKN, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNSX2 ( SI, SE, D, CKN, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNSX4 ( SI, SE, D, CKN, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNSXL ( SI, SE, D, CKN, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNX1 ( SI, SE, D, CKN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNX2 ( SI, SE, D, CKN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNX4 ( SI, SE, D, CKN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFNXL ( SI, SE, D, CKN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CKN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFRHQX1 ( SI, SE, D, CK, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule

module SDFFRHQX2 ( SI, SE, D, CK, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule

module SDFFRHQX4 ( SI, SE, D, CK, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule

module SDFFRHQXL ( SI, SE, D, CK, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;

endmodule

module SDFFRX1 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFRX2 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFRX4 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFRXL ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFSHQX1 ( SI, SE, D, CK, SN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule

module SDFFSHQX2 ( SI, SE, D, CK, SN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule

module SDFFSHQX4 ( SI, SE, D, CK, SN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule

module SDFFSHQXL ( SI, SE, D, CK, SN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;

endmodule

module SDFFSRHQX1 ( SI, SE, D, CK, SN, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule

module SDFFSRHQX2 ( SI, SE, D, CK, SN, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule

module SDFFSRHQX4 ( SI, SE, D, CK, SN, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule

module SDFFSRHQXL ( SI, SE, D, CK, SN, RN, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;

endmodule

module SDFFSRX1 ( SI, SE, D, CK, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFSRX2 ( SI, SE, D, CK, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFSRX4 ( SI, SE, D, CK, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFSRXL ( SI, SE, D, CK, SN, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFSX1 ( SI, SE, D, CK, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFSX2 ( SI, SE, D, CK, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFSX4 ( SI, SE, D, CK, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFSXL ( SI, SE, D, CK, SN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFTRX1 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFTRX2 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFTRX4 ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFTRXL ( SI, SE, D, CK, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SDFFX1 ( SI, SE, D, CK, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module SDFFX2 ( SI, SE, D, CK, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module SDFFX4 ( SI, SE, D, CK, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module SDFFXL ( SI, SE, D, CK, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    output		Q ;
    output		QN ;

endmodule

module SEDFFHQX1 ( SI, SE, D, CK, E, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;

endmodule

module SEDFFHQX2 ( SI, SE, D, CK, E, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;

endmodule

module SEDFFHQX4 ( SI, SE, D, CK, E, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;

endmodule

module SEDFFHQXL ( SI, SE, D, CK, E, Q);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;

endmodule

module SEDFFTRX1 ( SI, SE, D, CK, E, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SEDFFTRX2 ( SI, SE, D, CK, E, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SEDFFTRX4 ( SI, SE, D, CK, E, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SEDFFTRXL ( SI, SE, D, CK, E, RN, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module SEDFFX1 ( SI, SE, D, CK, E, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule

module SEDFFX2 ( SI, SE, D, CK, E, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule

module SEDFFX4 ( SI, SE, D, CK, E, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule

module SEDFFXL ( SI, SE, D, CK, E, Q, QN);
    input		SI ;
    input		SE ;
    input		D ;
    input		CK ;
    input		E ;
    output		Q ;
    output		QN ;

endmodule

module TBUFIX1 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFIX12 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFIX16 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFIX2 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFIX20 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFIX3 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFIX4 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFIX8 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFIXL ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFX1 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFX12 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFX16 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFX2 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFX20 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFX3 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFX4 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFX8 ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TBUFXL ( A, OE, Y);
    input		A ;
    input		OE ;
    output		Y ;

endmodule

module TIEHI ( Y);
    output		Y ;

endmodule

module TIELO ( Y);
    output		Y ;

endmodule

module TLATNRX1 ( D, GN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNRX2 ( D, GN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNRX4 ( D, GN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNRXL ( D, GN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNSRX1 ( D, GN, SN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNSRX2 ( D, GN, SN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNSRX4 ( D, GN, SN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNSRXL ( D, GN, SN, RN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNSX1 ( D, GN, SN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNSX2 ( D, GN, SN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNSX4 ( D, GN, SN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNSXL ( D, GN, SN, Q, QN);
    input		D ;
    input		GN ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNX1 ( D, GN, Q, QN);
    input		D ;
    input		GN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNX2 ( D, GN, Q, QN);
    input		D ;
    input		GN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNX4 ( D, GN, Q, QN);
    input		D ;
    input		GN ;
    output		Q ;
    output		QN ;

endmodule

module TLATNXL ( D, GN, Q, QN);
    input		D ;
    input		GN ;
    output		Q ;
    output		QN ;

endmodule

module TLATRX1 ( D, G, RN, Q, QN);
    input		D ;
    input		G ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATRX2 ( D, G, RN, Q, QN);
    input		D ;
    input		G ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATRX4 ( D, G, RN, Q, QN);
    input		D ;
    input		G ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATRXL ( D, G, RN, Q, QN);
    input		D ;
    input		G ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATSRX1 ( D, G, SN, RN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATSRX2 ( D, G, SN, RN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATSRX4 ( D, G, SN, RN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATSRXL ( D, G, SN, RN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    input		RN ;
    output		Q ;
    output		QN ;

endmodule

module TLATSX1 ( D, G, SN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module TLATSX2 ( D, G, SN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module TLATSX4 ( D, G, SN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module TLATSXL ( D, G, SN, Q, QN);
    input		D ;
    input		G ;
    input		SN ;
    output		Q ;
    output		QN ;

endmodule

module TLATX1 ( D, G, Q, QN);
    input		D ;
    input		G ;
    output		Q ;
    output		QN ;

endmodule

module TLATX2 ( D, G, Q, QN);
    input		D ;
    input		G ;
    output		Q ;
    output		QN ;

endmodule

module TLATX4 ( D, G, Q, QN);
    input		D ;
    input		G ;
    output		Q ;
    output		QN ;

endmodule

module TLATXL ( D, G, Q, QN);
    input		D ;
    input		G ;
    output		Q ;
    output		QN ;

endmodule

module TTLATX1 ( D, G, OE, Q);
    input		D ;
    input		G ;
    input		OE ;
    output		Q ;

endmodule

module TTLATX2 ( D, G, OE, Q);
    input		D ;
    input		G ;
    input		OE ;
    output		Q ;

endmodule

module TTLATX4 ( D, G, OE, Q);
    input		D ;
    input		G ;
    input		OE ;
    output		Q ;

endmodule

module TTLATXL ( D, G, OE, Q);
    input		D ;
    input		G ;
    input		OE ;
    output		Q ;

endmodule

module XNOR2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module XNOR2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module XNOR2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module XNOR2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module XNOR3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module XNOR3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module XOR2X1 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module XOR2X2 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module XOR2X4 ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module XOR2XL ( A, B, Y);
    input		A ;
    input		B ;
    output		Y ;

endmodule

module XOR3X2 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module XOR3X4 ( A, B, C, Y);
    input		A ;
    input		B ;
    input		C ;
    output		Y ;

endmodule

module PDB04DGZ ( I, OEN, PAD, C);
    input		I ;
    input		OEN ;
    inout		PAD ;
    output		C ;

endmodule

module PDIDGZ ( PAD, C);
    input		PAD ;
    output		C ;

endmodule

module PDO04CDG ( I, PAD);
    input		I ;
    output		PAD ;

endmodule

module PVDD1DGZ ( );

endmodule

module PVSS1DGZ ( );

endmodule

module pllclk ( refclk, ibias, reset, clk1x, clk2x, vcop, vcom);
    input		refclk ;
    input		ibias ;
    input		reset ;
    output		clk1x ;
    output		clk2x ;
    output		vcop ;
    output		vcom ;

endmodule

module ram_128x16A ( CEN, OEN, WEN, CLK, Q, A, D);
    input		CEN ;
    input		OEN ;
    input		WEN ;
    input		CLK ;
    output  [15:0]  Q ;
    input  [6:0]  A ;
    input  [15:0]  D ;

endmodule

module ram_256x16A ( CEN, OEN, WEN, CLK, Q, A, D);
    input		CEN ;
    input		OEN ;
    input		WEN ;
    input		CLK ;
    output  [15:0]  Q ;
    input  [7:0]  A ;
    input  [15:0]  D ;

endmodule

module rom_512x16A ( CEN, CLK, Q, A);
    input		CEN ;
    input		CLK ;
    output  [15:0]  Q ;
    input  [8:0]  A ;

endmodule

module PCORNERDG ( );

endmodule
